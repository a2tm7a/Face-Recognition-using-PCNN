--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

library work;
use work.arraypack.all;

package inputs is

procedure get_input(variable x_2D  : out x_array_2D;
						 variable w_2D  : out w_array_2D;
						 variable yp_2D  : out yp_array_2D);

procedure calculate_y(variable x_1D : in x_array_1D;
							 variable w_2D : in w_array_2D;
							 variable y_1D : out y_array_1D);

procedure distance(variable y_1D : in y_array_1D;
						 variable yp_2D : in yp_array_2D;
						 variable index : out integer;
						 variable minNorm : out integer);
							
end inputs;

package body inputs is
	
	procedure get_input(variable x_2D  : out x_array_2D;
								variable w_2D  : out w_array_2D;
								variable yp_2D  : out yp_array_2D) IS
		begin
			x_2D := ((8,7,6,6,5,5,6,7,9,11,9,9,9,10,7,8,9,6,6,7,6,6,5,5,5,5,4,4,5,4,5,5,6,5,5,5,5,4,4,8,12,13,13,12,10,10,10,6,8,7,8,6,7,7,4,4,4,5,5,6,6,4,3,4,4,2,3,4,4,4,6,12,13,13,12,14,11,10,10,8,8,8,8,8,7,6,5,6,6,7,5,4,4,4,4,4,4,2,1,2,4,6,9,12,13,14,14,12,12,8,8,8,8,10,9,8,7,8,6,5,5,7,5,3,3,3,3,4,5,2,2,3,4,7,11,12,13,14,13,13,12,9,9,7,7,10,12,11,9,7,6,5,5,5,4,3,1,2,3,3,3,2,2,3,4,6,10,13,14,14,14,14,12,12,7,8,8,9,10,10,11,8,7,6,5,4,3,3,3,1,2,3,3,2,2,2,3,5,10,13,14,15,15,15,15,12,9,8,9,11,11,12,12,11,9,8,7,5,2,2,1,3,2,3,4,2,1,1,2,5,11,14,15,16,15,15,14,14,11,8,9,11,13,15,12,11,10,9,7,6,2,1,1,1,2,2,1,1,0,2,3,6,13,16,17,16,15,14,13,13,12,10,8,11,13,13,12,12,12,10,10,7,2,1,1,1,3,0,2,0,1,3,1,9,13,15,14,13,11,9,11,10,11,10,10,11,12,12,13,14,15,13,11,8,4,0,1,1,2,1,2,2,2,2,1,11,12,9,7,4,3,3,4,6,7,8,10,9,7,6,6,5,7,9,10,9,5,0,1,1,1,2,3,2,3,0,3,12,8,6,5,7,6,3,2,3,5,13,13,6,3,2,1,2,3,4,5,9,6,0,1,0,1,3,6,3,3,0,9,12,9,6,7,8,8,4,2,2,5,19,19,7,2,1,2,5,4,4,3,5,8,2,0,0,1,2,13,7,4,1,11,13,12,9,5,5,4,5,6,7,11,19,18,10,5,3,2,2,3,5,4,6,8,5,0,0,0,3,19,17,5,2,13,14,14,14,12,11,12,13,12,15,12,19,18,10,13,9,7,7,6,6,8,9,10,8,0,0,1,3,19,19,7,5,13,15,17,18,18,19,19,19,18,15,12,19,16,10,13,16,17,16,14,13,13,13,12,9,1,1,2,3,19,19,8,8,12,14,17,19,19,19,19,19,17,14,14,18,16,11,12,15,19,19,19,18,17,14,13,10,3,2,3,6,19,19,8,10,12,12,15,16,19,19,19,19,13,11,14,19,19,12,10,13,19,19,19,18,16,14,12,10,7,2,7,19,19,19,11,10,12,12,14,15,18,19,19,18,10,14,13,16,15,12,13,10,17,19,19,17,14,12,10,10,9,1,17,18,19,19,11,12,12,12,13,14,15,17,17,15,9,7,6,8,6,5,9,9,15,16,16,14,12,11,10,9,9,2,18,19,19,19,12,13,11,12,12,12,13,14,14,15,12,2,1,3,2,0,1,11,14,13,13,12,11,10,10,9,9,6,16,19,19,19,19,13,11,11,11,11,13,14,16,13,10,10,8,3,3,8,8,10,13,13,12,10,9,9,9,9,9,7,19,19,19,19,19,8,11,10,11,11,14,14,15,12,11,12,10,8,7,11,10,10,11,13,12,10,10,9,9,9,9,14,16,19,19,19,19,3,11,10,10,11,14,13,12,11,11,8,10,15,15,9,10,10,9,11,12,11,10,8,8,9,5,19,19,17,19,19,19,16,11,10,10,12,14,14,6,4,3,2,3,2,2,3,4,4,5,8,11,12,10,8,8,8,17,16,19,19,19,19,19,18,15,10,10,12,14,12,9,9,7,9,10,10,8,8,7,4,3,5,9,11,10,8,8,8,19,19,18,19,19,19,19,19,19,10,10,11,12,11,12,13,12,10,6,5,4,6,8,10,11,11,9,10,9,8,8,9,19,19,19,19,19,19,19,19,18,9,10,10,10,11,10,11,10,8,7,6,5,7,8,9,10,10,9,8,8,8,7,19,19,19,19,19,19,19,19,19,19,12,9,10,9,9,11,10,9,9,7,6,6,7,8,8,8,8,9,8,8,8,7,19,19,19,18,19,19,19,19,19,19,14,9,9,9,10,12,13,14,17,18,18,17,16,12,10,10,9,8,8,8,7,19,19,19,19,19,19,19,19,19,19,19,14,10,7,8,8,12,14,15,18,18,14,16,19,16,15,12,9,7,7,6,17,19,19,18,19,19,19,19,19,19,19,19,14,11,7,6,7,9,11,12,12,12,11,12,13,12,12,10,8,6,5,6,18,19,19,19,19,19,19),(19,1,0,0,0,2,8,10,11,11,12,13,15,14,15,14,14,16,15,15,13,11,10,8,8,7,4,0,0,0,0,0,8,1,0,0,0,6,9,10,11,11,12,14,16,15,14,14,14,15,16,16,14,11,10,8,8,7,6,2,0,0,0,0,2,0,0,0,1,7,10,10,10,11,12,13,15,14,15,14,13,14,14,15,13,10,10,8,8,7,6,4,0,0,0,0,1,1,0,0,2,7,9,10,10,11,11,12,14,13,13,13,12,13,12,13,11,9,9,9,7,7,7,5,1,0,0,0,0,1,0,0,3,8,9,10,10,11,11,12,13,13,14,13,13,13,13,12,11,9,9,8,7,7,6,5,2,0,0,0,0,1,0,0,3,8,9,9,10,11,12,13,14,14,13,13,13,13,13,14,12,10,9,9,8,7,6,5,2,0,0,0,1,1,1,0,3,8,8,9,10,11,12,13,14,15,14,14,14,13,13,13,11,10,10,8,8,7,6,5,1,0,0,0,0,0,1,0,4,9,9,10,9,11,12,13,14,13,13,13,14,15,13,12,12,11,10,9,8,7,6,6,1,0,0,0,0,0,0,0,6,9,9,9,6,7,8,10,11,11,11,11,12,12,11,10,11,9,8,8,7,7,6,6,1,0,0,0,2,0,0,0,8,8,7,3,2,2,2,2,5,8,10,10,11,10,10,8,7,5,4,3,3,4,6,6,1,0,0,0,13,1,0,1,9,8,4,3,3,2,1,1,1,2,5,8,10,7,5,3,2,1,1,1,1,1,3,6,3,0,0,2,18,6,0,1,10,7,4,4,4,4,3,1,1,2,4,9,9,6,3,2,1,1,1,1,2,2,2,5,4,0,0,8,5,4,3,2,10,8,5,4,3,4,3,2,1,1,5,12,11,8,3,0,0,1,2,2,2,2,3,5,5,0,3,8,4,7,5,3,10,9,7,6,3,1,0,1,3,4,5,12,14,9,2,1,0,1,2,2,2,2,3,5,6,0,4,3,6,8,6,5,10,9,9,8,7,5,6,6,6,6,7,12,14,9,4,3,2,1,1,1,3,5,5,6,6,1,4,2,7,9,5,9,9,10,11,12,13,12,11,8,11,9,9,13,14,8,5,6,5,6,6,5,6,7,7,6,6,4,5,3,7,6,5,10,10,10,10,10,12,12,12,12,11,9,9,13,12,8,6,6,8,7,7,8,8,7,7,6,6,2,5,4,8,6,8,9,9,9,9,9,10,12,13,12,10,8,10,12,12,8,6,6,9,9,9,9,8,7,6,6,6,3,4,4,7,10,9,8,9,8,8,9,11,12,12,11,9,9,10,14,13,8,6,5,8,9,9,9,7,6,5,6,6,6,5,5,11,9,9,8,9,8,7,7,10,11,12,10,8,8,7,9,8,7,6,6,7,8,9,8,6,6,5,5,5,6,7,5,19,11,11,8,8,8,8,8,9,10,9,8,6,4,3,5,4,4,3,5,5,7,7,7,6,5,5,5,6,6,4,8,19,10,8,16,8,7,7,7,8,9,8,9,8,2,1,2,1,1,1,5,6,6,7,6,5,5,5,5,6,7,8,17,19,19,19,19,8,7,7,7,7,8,9,9,6,2,1,1,0,1,1,5,6,7,6,6,5,5,5,5,12,5,8,16,19,19,19,19,8,7,7,7,7,8,4,4,3,1,1,1,1,1,1,2,4,4,5,5,5,5,5,6,15,16,14,16,19,19,19,19,9,7,7,7,7,5,1,2,1,1,1,1,0,1,1,1,1,1,3,5,4,4,5,10,15,15,15,17,19,19,19,18,9,7,7,7,6,3,1,1,1,1,2,1,0,1,1,1,1,0,1,4,4,5,5,15,15,16,15,15,19,19,19,19,13,7,7,7,7,3,1,1,2,1,1,1,0,0,0,0,0,0,1,4,4,4,5,14,15,17,16,14,19,19,19,19,19,7,7,6,6,5,4,4,5,4,5,4,4,4,3,3,3,2,3,4,4,4,6,17,16,16,16,15,19,19,19,19,19,10,6,6,6,4,4,4,4,3,2,1,1,2,2,3,3,3,3,4,4,4,13,17,16,16,15,16,19,19,19,19,19,19,6,6,6,5,5,4,5,4,2,2,2,2,3,4,3,3,4,4,4,5,17,19,18,15,17,15,19,19,19,19,19,18,7,6,6,6,6,6,7,8,9,9,9,7,7,5,4,4,4,4,4,6,18,16,18,15,16,15,19,19,19,19,19,9,8,5,6,6,6,6,7,8,10,8,7,7,6,5,5,4,4,4,3,6,16,18,17,16,16,14),(2,2,1,1,1,0,0,0,2,7,12,15,13,13,11,10,7,4,2,2,1,1,0,0,0,1,1,1,0,0,0,1,1,1,1,1,0,0,1,2,7,13,15,17,17,16,14,13,11,8,5,4,2,1,0,0,0,0,0,1,0,0,0,0,1,0,0,1,0,0,1,8,13,15,17,18,17,16,15,13,12,10,8,6,3,2,1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,3,11,14,15,16,16,17,16,16,14,13,11,10,8,4,2,1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,6,11,14,16,15,16,16,17,17,15,15,14,10,9,6,3,1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,1,8,12,14,16,17,18,18,18,18,17,17,16,14,11,9,4,3,1,1,0,0,0,0,0,0,0,0,0,0,0,0,2,8,12,14,17,17,18,19,19,18,18,18,17,16,13,11,8,4,3,1,1,1,1,0,0,0,0,1,0,0,0,0,5,9,12,15,17,17,17,18,18,18,18,19,18,17,16,13,11,5,5,3,1,0,0,0,0,0,0,1,0,0,0,2,7,9,13,14,15,15,14,13,14,15,15,17,16,14,13,13,11,8,5,5,3,2,2,0,0,0,0,0,0,0,0,4,9,11,8,7,5,6,6,7,9,11,12,12,12,8,6,5,4,3,3,4,5,4,2,1,0,0,0,1,0,0,0,6,10,8,3,2,1,1,1,1,3,8,11,12,8,3,1,1,1,1,2,2,4,5,4,2,0,0,0,1,0,1,2,9,9,5,6,7,8,6,4,3,3,7,14,14,6,3,3,3,4,5,6,5,4,5,6,4,0,0,0,2,1,0,4,11,9,8,8,9,13,13,7,3,3,7,16,16,7,2,3,5,9,11,9,7,7,6,7,7,1,0,0,3,2,1,6,11,9,8,7,8,7,7,4,2,5,7,17,18,7,3,2,4,8,8,7,6,6,7,8,9,3,0,0,7,4,1,7,11,10,9,7,2,2,2,2,6,9,9,18,18,8,9,6,2,2,2,3,4,7,8,9,9,3,0,1,17,6,1,8,12,11,11,10,5,4,4,6,11,11,10,19,18,8,10,12,7,4,4,5,8,9,9,9,9,3,0,1,19,9,4,9,12,12,13,13,13,12,11,13,13,10,11,19,16,8,9,13,12,10,9,10,11,12,11,9,9,2,0,2,19,11,6,8,12,11,12,13,15,16,15,13,11,9,9,17,15,9,8,9,12,12,13,13,13,12,11,9,9,2,2,4,19,13,10,6,11,10,11,13,14,16,14,14,10,8,9,16,15,9,7,9,12,13,14,13,12,10,8,8,9,5,5,7,19,19,11,8,11,10,10,11,12,13,13,12,7,9,11,16,15,9,8,6,10,12,12,12,10,8,7,7,8,5,7,8,19,19,15,8,10,9,9,9,10,11,11,10,9,11,12,17,17,10,10,8,9,11,11,9,8,7,7,7,7,5,4,9,19,19,19,14,9,9,9,8,9,10,10,11,7,7,11,12,13,9,5,6,9,10,9,8,7,7,7,7,7,7,9,19,19,19,19,19,11,9,8,8,9,10,12,11,8,3,3,5,4,2,2,8,9,10,8,7,7,7,7,7,7,18,19,19,19,19,19,19,12,9,8,8,9,10,11,10,9,6,3,1,2,2,5,8,10,10,8,8,7,7,7,7,8,18,19,19,19,19,19,19,16,9,8,9,10,9,8,6,7,6,6,4,3,5,5,6,7,8,8,8,8,7,7,7,11,19,19,19,19,19,19,19,19,9,8,9,9,6,6,5,5,4,4,5,3,4,5,7,7,6,8,8,8,7,7,7,15,19,19,19,19,19,19,19,19,9,8,8,9,6,3,2,2,2,3,2,3,4,2,1,2,6,7,8,8,7,7,6,19,19,19,19,19,19,19,19,19,14,7,8,8,7,7,7,6,8,11,10,8,7,6,6,6,5,7,8,7,6,6,7,19,19,19,19,19,19,19,19,19,19,7,7,8,7,7,7,6,6,6,6,5,5,5,6,7,6,7,7,7,5,6,9,19,19,19,19,19,19,19,19,19,19,12,6,7,6,6,7,6,4,2,1,2,3,5,6,7,6,6,6,6,4,4,14,19,19,19,19,19,19,19,19,19,19,14,4,6,6,6,7,6,6,5,3,4,5,6,7,6,5,6,5,4,3,6,8,19,19,19,19,19,19,19,19,19,19,7,8,3,4,5,8,9,9,11,8,9,10,9,8,7,4,6,4,2,3,6,3,19,19,19,19),(19,19,12,2,2,1,1,1,1,1,1,0,0,0,1,1,2,3,5,5,5,4,3,2,1,0,0,0,0,0,0,1,19,19,1,1,0,0,1,0,1,1,0,0,1,2,2,4,6,8,9,9,8,7,6,3,1,0,0,0,0,0,0,0,19,10,1,1,0,0,1,1,0,0,0,1,2,4,5,7,8,9,9,9,8,7,6,4,2,1,0,0,0,0,0,0,19,1,1,0,0,0,0,1,0,0,1,2,4,5,6,8,9,9,9,9,8,7,6,5,3,2,0,0,0,0,0,0,17,1,0,0,0,0,0,0,0,0,2,3,6,6,7,8,9,9,9,9,9,7,6,5,4,3,0,0,0,0,0,0,4,1,0,0,0,0,0,0,0,1,4,6,7,8,9,9,10,10,10,10,9,8,7,6,5,4,1,0,0,0,0,0,1,0,0,0,0,0,0,0,2,5,7,10,9,10,11,10,12,11,10,11,10,9,7,6,5,4,1,1,0,0,0,0,1,0,0,0,0,0,1,2,3,9,10,10,9,10,11,11,11,12,10,10,10,9,8,7,6,4,1,0,0,0,0,0,1,0,0,0,0,3,1,2,3,3,5,8,8,9,9,10,10,10,9,9,9,9,8,8,6,5,1,0,0,0,0,0,1,0,0,1,5,6,2,3,3,4,4,4,4,6,8,9,9,8,7,6,4,3,3,3,3,5,2,0,0,0,0,0,1,1,0,6,8,7,5,6,8,10,9,6,5,4,7,10,9,7,4,3,3,3,4,3,2,5,3,1,0,0,0,0,1,1,0,8,8,7,6,6,7,10,10,8,7,7,8,10,9,7,5,6,6,9,8,6,4,5,5,2,0,0,0,1,2,1,1,10,9,7,4,3,4,6,4,4,7,7,9,12,11,7,6,6,7,9,8,6,5,5,6,5,0,0,0,8,3,1,4,9,9,9,9,6,4,3,4,6,8,9,9,13,12,8,7,7,1,3,4,3,3,4,6,7,2,0,1,17,4,2,7,10,10,11,10,10,9,9,10,10,11,9,9,13,11,8,8,8,8,5,3,4,6,6,7,7,4,0,1,15,8,5,9,10,11,11,11,11,11,10,11,12,11,9,10,13,12,8,8,10,10,8,8,8,8,8,8,7,6,1,1,16,9,3,10,10,10,11,12,12,12,12,13,12,10,9,10,12,11,8,8,10,11,10,9,10,9,9,8,7,7,2,2,19,10,6,10,9,9,10,11,14,14,13,12,11,9,8,10,12,12,9,7,8,10,11,10,10,10,9,8,8,7,3,4,15,10,9,9,8,9,9,11,13,14,13,12,9,7,9,12,14,13,9,7,7,10,11,11,10,10,8,8,7,7,5,6,15,12,10,9,8,9,9,9,10,12,12,11,9,10,9,7,9,8,7,9,6,9,10,10,9,9,7,7,7,7,7,15,17,19,11,9,8,8,8,9,10,10,11,11,7,7,2,4,4,4,3,7,6,9,9,10,9,7,6,6,7,7,5,19,16,18,10,10,8,8,8,9,9,9,11,11,8,3,3,3,2,2,1,3,6,9,9,8,7,7,6,6,7,7,8,19,17,19,19,10,8,8,9,9,9,9,10,11,9,9,7,8,6,8,7,6,8,8,9,7,7,6,6,5,6,8,18,19,17,19,17,12,8,8,9,9,9,9,9,10,10,9,10,9,9,10,9,8,8,9,8,7,7,6,6,6,6,13,19,15,19,17,19,18,8,9,9,9,8,7,7,7,8,8,5,7,8,8,8,8,7,8,7,6,7,6,6,6,9,19,19,18,17,19,17,19,8,8,9,8,7,7,6,3,3,2,2,2,3,2,2,4,6,5,6,6,6,6,6,6,15,17,18,18,15,19,19,19,8,8,8,8,7,7,5,4,2,3,3,1,1,1,1,1,1,4,5,6,6,6,6,6,17,15,16,16,16,19,19,19,16,7,7,7,7,6,6,7,5,5,8,8,9,8,4,3,5,4,5,6,6,6,5,11,18,15,19,15,19,19,17,15,15,6,6,6,6,6,6,6,5,3,3,4,4,3,3,4,5,5,5,5,5,5,5,14,19,19,16,19,19,17,18,19,19,14,5,5,5,5,5,5,5,4,2,2,2,2,3,4,5,5,4,4,5,4,14,16,19,16,19,15,17,19,18,18,18,16,5,4,5,6,5,5,5,5,6,4,3,4,5,5,5,4,4,4,4,4,17,15,16,16,19,19,19,19,18,19,19,18,6,3,4,5,6,6,6,6,7,6,6,6,6,5,5,5,4,3,3,5,12,15,18,19,18,19,17),(19,19,19,19,7,5,5,11,13,13,13,13,14,15,14,14,14,15,14,13,12,11,12,12,12,11,7,18,19,19,19,19,19,19,19,7,6,4,11,12,12,13,13,13,15,15,15,16,16,14,14,13,13,12,11,11,11,11,11,11,19,19,19,19,19,19,11,7,5,6,11,12,12,12,13,14,15,16,16,17,17,16,15,14,15,13,11,10,10,10,10,8,10,18,19,19,19,16,6,9,5,9,11,11,11,12,13,14,15,16,15,16,16,15,15,15,14,11,10,10,8,9,9,9,6,10,19,19,19,10,7,7,6,10,10,11,11,12,11,13,15,15,15,15,15,15,14,15,14,11,10,10,10,9,8,8,5,7,8,19,19,7,6,7,8,10,9,11,11,11,12,14,14,15,15,15,16,15,14,14,13,12,10,10,10,8,8,8,6,6,9,19,19,7,6,8,8,9,9,10,11,11,13,14,15,15,16,15,15,13,14,14,14,11,11,10,10,7,7,7,6,6,8,9,19,7,5,8,8,9,8,10,12,12,12,13,12,14,15,15,14,14,12,13,13,12,11,10,9,7,7,7,6,5,6,8,19,6,7,9,9,8,8,9,10,11,11,11,10,10,12,13,11,12,8,9,7,8,8,7,8,7,6,7,7,6,6,7,19,7,6,8,7,8,8,8,5,5,4,3,3,4,9,12,9,8,4,2,2,3,3,4,4,6,7,6,7,6,5,7,19,8,9,8,7,8,7,3,3,2,1,1,1,2,5,11,9,4,2,1,1,1,2,3,3,5,6,6,5,6,6,7,19,10,8,8,8,8,5,3,5,6,4,3,2,2,6,13,11,3,1,1,2,4,5,3,4,5,6,6,5,6,6,7,19,13,9,9,8,9,4,4,6,7,10,6,2,2,6,10,10,3,1,2,5,8,6,5,3,4,6,7,5,5,6,9,19,15,8,8,9,9,7,6,5,5,6,4,3,4,6,10,9,5,4,1,3,5,4,5,4,5,6,7,7,4,5,8,19,19,9,10,10,9,7,6,3,2,1,2,5,7,7,10,9,6,7,5,2,1,1,3,5,6,6,8,8,4,3,12,19,13,11,13,11,9,10,10,8,6,6,5,8,8,7,11,10,6,8,9,7,5,6,7,8,8,8,8,8,10,7,7,19,5,9,12,10,10,14,12,11,11,10,10,10,7,8,11,12,7,7,10,11,7,9,11,10,11,9,8,8,10,6,2,19,5,9,10,10,9,12,13,11,11,11,12,8,7,7,11,11,8,6,9,10,9,8,8,9,10,7,7,7,9,5,6,19,8,7,9,9,8,8,9,9,9,11,11,7,8,8,10,9,7,7,7,10,8,8,8,8,7,6,6,6,8,4,6,19,11,5,10,9,7,6,7,8,10,10,10,6,6,6,5,4,4,4,4,8,9,7,7,5,5,6,6,7,7,2,4,19,10,6,9,10,7,6,6,8,9,10,7,5,3,0,4,4,0,2,5,5,8,7,6,5,5,6,7,7,6,3,4,19,13,7,9,10,8,7,7,8,9,8,7,7,2,3,2,1,4,4,6,6,6,7,7,5,6,6,7,6,6,5,6,19,19,9,9,10,8,7,7,8,8,5,7,8,7,6,5,4,6,6,7,6,3,7,7,6,5,6,6,6,4,7,5,19,19,11,9,9,8,8,9,8,7,6,7,6,6,6,5,6,6,6,6,6,5,5,6,5,6,6,6,6,5,5,10,19,19,13,7,9,8,7,7,8,6,6,6,6,6,6,6,7,6,5,5,6,5,4,6,6,6,5,6,6,7,8,17,19,19,19,7,8,8,7,7,7,5,6,6,5,5,4,5,5,4,4,5,5,5,4,5,5,6,6,6,6,7,14,17,19,19,19,19,10,8,8,7,7,4,5,5,3,2,2,1,2,2,2,2,3,4,3,5,5,6,6,5,19,17,19,19,19,19,19,19,18,8,8,7,7,5,5,1,1,2,4,4,5,4,3,3,2,4,4,6,5,6,6,5,19,19,17,18,19,19,19,19,19,8,8,8,8,6,5,6,7,6,5,4,4,5,5,5,4,4,5,6,5,6,5,6,18,19,19,18,19,19,19,19,19,12,8,8,7,6,5,6,5,4,3,3,3,3,3,4,5,5,5,5,5,6,4,11,19,19,18,18,19,19,19,19,19,15,7,8,7,6,5,5,4,3,2,2,2,3,4,4,5,5,5,5,6,5,5,12,19,19,19,19,19,19,19,19,19,8,7,8,7,6,6,5,5,4,10,10,10,8,5,6,5,5,5,5,6,5,5,7,19,17,19,19),(17,0,0,0,0,0,0,0,0,0,1,2,4,5,6,7,6,6,6,7,7,7,6,6,5,3,0,1,1,1,1,2,5,0,0,0,0,0,0,0,2,4,8,10,10,10,11,11,11,11,11,11,9,9,8,7,7,5,2,0,0,1,1,1,0,0,0,0,0,0,2,4,7,9,11,13,12,12,12,12,11,12,12,12,11,10,9,8,7,6,3,0,0,0,1,1,0,0,0,0,0,3,6,7,8,9,11,12,12,12,12,12,12,12,12,13,13,11,9,8,7,6,5,1,0,0,0,1,0,0,0,0,0,4,6,8,9,9,11,12,12,12,12,12,12,12,12,12,12,11,9,8,7,6,5,3,0,0,0,0,0,0,0,0,2,5,6,8,9,9,10,12,12,12,12,12,12,12,13,13,12,11,10,9,7,6,6,4,1,0,0,0,0,0,0,0,3,5,6,7,9,10,11,12,13,12,12,12,14,13,13,14,14,12,11,9,7,6,6,5,2,0,0,0,0,0,0,1,3,5,6,7,9,11,12,14,14,13,13,13,14,14,14,14,12,10,9,7,7,6,6,5,3,0,0,0,0,0,0,1,4,5,6,5,6,6,6,6,8,10,11,11,11,11,9,4,2,2,3,4,5,6,6,5,5,1,0,0,0,0,0,2,5,5,4,3,3,1,1,1,3,6,7,8,8,7,4,3,2,2,2,3,4,5,6,6,5,3,0,0,0,0,0,3,5,5,4,4,3,3,3,3,3,3,5,8,9,6,3,3,6,9,10,7,5,4,6,6,6,4,0,0,0,0,0,4,5,5,4,4,7,10,8,7,4,4,7,11,12,8,4,5,7,9,9,7,6,5,5,6,7,5,0,0,0,0,0,4,5,5,4,5,6,6,4,3,4,5,8,12,13,8,6,4,1,2,2,3,4,5,6,7,7,6,1,0,0,0,0,5,6,5,4,3,1,0,1,3,4,8,7,11,12,8,7,7,4,4,4,4,4,5,7,8,7,7,1,0,0,0,0,5,6,6,3,3,4,4,4,3,6,8,7,12,13,8,8,9,7,5,5,6,7,9,11,9,8,7,2,1,0,0,0,6,7,8,8,8,7,6,8,9,8,9,7,12,13,8,9,8,10,11,11,11,12,11,11,10,8,7,4,0,0,0,0,6,8,9,10,10,12,12,12,11,8,9,8,12,12,8,7,7,9,11,12,12,12,11,10,9,8,7,7,3,2,0,1,7,8,9,9,11,12,11,11,11,8,6,8,14,15,9,7,5,9,11,12,11,11,10,9,8,7,7,7,3,3,2,3,7,6,8,9,10,11,11,12,10,7,9,7,8,8,7,9,9,7,10,12,11,12,10,8,7,6,6,7,1,5,3,2,6,6,7,8,9,10,10,9,8,6,5,2,4,4,4,4,6,6,8,10,11,10,9,7,6,6,6,7,5,7,3,6,6,5,6,7,8,8,8,7,6,4,1,1,2,2,1,1,2,6,7,8,9,8,7,6,5,6,6,7,7,7,5,6,6,5,5,6,7,7,7,6,7,7,6,7,6,5,7,7,7,8,9,7,7,7,7,6,6,6,6,7,8,6,6,7,6,6,5,5,6,6,6,7,8,8,7,8,9,8,9,8,8,9,9,9,6,7,6,5,6,6,6,7,7,7,5,7,6,5,6,5,5,5,6,7,7,7,8,9,10,10,11,9,8,7,7,8,8,6,6,6,6,6,7,7,8,15,8,8,7,6,6,6,6,6,8,6,5,5,4,3,3,2,3,2,2,4,4,6,7,6,6,6,6,6,7,5,7,17,14,7,6,6,6,6,6,6,7,5,1,0,1,1,1,1,2,2,3,1,3,5,7,7,6,6,6,6,7,0,8,14,13,8,0,6,6,6,6,6,7,5,6,4,3,4,6,6,5,3,4,5,7,7,7,7,6,6,5,6,5,2,14,16,15,14,5,5,6,6,6,6,6,7,7,6,4,3,2,2,2,3,5,7,8,7,6,6,6,5,5,5,1,13,18,16,17,19,15,5,5,5,5,5,5,7,8,7,6,6,5,5,5,6,7,8,7,6,5,5,5,5,5,4,7,14,15,15,14,16,13,6,4,4,4,5,5,7,7,8,8,9,9,10,10,9,8,8,7,6,5,5,5,4,4,4,15,14,17,14,15,19,15,15,9,4,4,4,5,4,8,8,10,11,11,11,11,11,11,9,8,6,5,5,4,3,5,14,17,14,14,14,15,14,14,17,14,13,3,4,4,5,6,8,8,9,8,9,8,8,7,6,6,5,4,3,3,3,6,15,14,16,15),(1,1,1,1,1,1,2,2,2,2,2,3,4,4,5,5,4,5,6,6,8,8,5,3,2,2,2,1,1,1,1,1,1,1,1,1,1,2,3,2,3,3,4,5,7,7,7,7,7,8,9,11,14,13,8,4,3,3,2,2,1,0,1,1,2,0,1,1,1,3,4,4,4,3,5,7,8,8,9,9,9,10,10,11,13,11,8,6,4,3,3,2,1,0,0,0,1,1,1,1,2,4,5,5,4,5,6,7,8,9,9,11,11,11,10,10,9,8,6,6,6,4,4,3,1,0,0,0,3,2,1,1,2,5,5,5,6,7,8,10,10,11,12,12,12,11,10,10,9,8,6,6,6,6,5,4,1,0,0,0,3,2,1,1,4,6,6,6,7,8,10,12,14,14,14,13,13,13,13,13,12,10,8,6,6,6,5,5,3,0,0,0,3,1,2,2,7,6,7,7,8,10,11,13,15,17,16,16,15,16,15,15,14,11,8,7,6,6,6,7,4,1,0,0,5,1,1,3,9,7,7,9,8,10,12,13,13,14,15,16,17,17,15,14,12,10,9,9,7,6,6,7,7,1,1,1,8,2,1,4,9,8,8,3,3,4,7,8,9,10,11,11,12,12,12,11,10,8,8,7,5,7,7,7,8,1,1,1,5,4,1,7,9,9,4,2,3,2,2,3,4,5,7,8,9,9,8,6,4,3,2,2,3,3,4,8,8,2,1,3,4,5,1,8,9,7,5,4,3,3,1,1,0,1,3,6,8,5,3,1,0,0,1,1,2,2,3,6,8,2,1,3,6,6,1,9,9,6,4,5,4,4,4,2,1,1,1,5,7,4,2,1,1,2,3,3,3,4,4,5,8,3,1,5,7,3,2,9,8,7,5,4,4,3,3,2,1,1,1,7,11,6,1,1,1,3,4,3,3,4,3,5,7,4,2,6,7,3,2,8,9,8,7,4,2,1,1,1,1,2,3,9,14,8,2,1,1,1,2,3,2,3,5,6,8,6,2,4,7,4,6,9,9,8,9,7,5,3,3,3,4,7,7,12,15,8,5,4,2,2,2,2,3,5,7,7,8,5,2,7,8,9,5,8,8,8,10,10,9,7,6,7,11,10,9,12,15,8,7,8,7,5,4,4,6,7,8,8,8,5,7,6,11,9,6,7,7,8,9,10,11,12,14,14,11,8,8,12,16,8,7,7,9,10,8,10,11,9,8,7,8,4,9,7,10,9,4,6,7,6,8,9,12,13,14,11,7,8,11,15,18,10,7,5,9,12,13,13,11,9,7,6,7,2,8,10,10,8,4,4,5,5,8,10,11,11,10,8,6,11,10,15,19,9,7,7,6,10,11,12,11,9,6,6,6,2,9,9,19,15,5,3,4,5,7,9,9,8,7,8,7,9,9,11,10,8,8,9,6,8,9,9,9,8,6,5,4,1,5,16,19,19,9,2,2,4,7,7,7,6,6,8,8,3,1,4,4,3,5,5,7,6,7,7,7,6,4,4,2,7,19,19,19,19,10,1,2,3,4,4,4,4,3,2,2,0,0,0,0,0,0,3,4,5,4,5,5,5,4,3,1,10,19,19,19,19,12,1,2,3,3,3,3,1,1,2,1,1,0,0,0,0,0,0,0,1,2,3,4,3,2,2,1,16,19,19,19,19,18,1,1,2,2,2,1,1,0,1,2,1,1,3,4,1,1,1,1,1,0,1,2,2,1,1,1,19,19,19,19,19,19,3,1,1,2,3,1,0,0,0,1,1,1,2,1,1,1,1,0,0,0,0,3,2,1,1,3,19,19,19,19,19,19,14,1,1,1,2,0,0,1,3,5,7,9,11,10,7,5,3,1,0,0,1,3,2,1,1,16,19,19,19,19,19,19,19,5,1,1,1,0,1,2,2,2,4,6,8,8,5,4,2,1,1,0,1,2,1,1,3,19,19,19,19,19,19,19,19,18,1,1,0,0,1,2,2,1,0,0,0,0,0,1,1,1,1,0,1,1,0,0,19,19,19,19,19,19,19,19,19,19,3,1,0,0,0,1,1,1,1,1,1,2,1,1,1,1,1,0,0,0,0,3,19,19,19,19,19,19,19,19,19,19,6,1,0,0,0,1,1,1,1,3,6,4,3,1,1,0,0,0,0,0,0,6,19,19,19,19,19,19,19,19,19,19,6,1,1,0,0,0,1,1,2,4,4,2,2,1,1,1,0,0,0,0,0,8,19,19,19,19,19,19,19,19,19,19,7,4,1,0,0,0,0,0,1,2,2,1,1,1,0,0,0,0,0,0,2,12,19,19,19,19,19),(19,19,1,1,1,0,0,0,0,1,1,6,12,13,14,15,15,15,15,14,12,10,6,4,3,2,1,1,1,1,4,19,19,15,1,1,0,0,0,1,1,5,13,15,15,16,15,15,16,16,15,15,13,12,8,4,5,4,1,0,0,1,2,19,19,2,0,0,0,1,7,1,8,12,14,16,15,16,15,15,15,15,15,14,13,12,10,7,5,4,3,1,0,0,1,2,19,1,0,0,0,8,4,9,10,11,14,15,15,15,15,15,15,15,14,13,12,11,10,10,7,5,6,1,0,0,0,1,19,0,0,0,6,6,9,10,10,12,13,15,16,15,15,15,14,14,14,14,13,12,11,10,9,7,3,3,0,0,0,1,16,0,0,5,8,7,9,10,11,12,13,16,16,16,16,15,16,16,15,15,14,13,11,10,10,8,8,3,1,0,0,0,12,0,1,5,8,8,9,10,11,13,15,15,16,16,16,16,16,16,16,15,15,14,12,10,9,8,9,7,2,0,0,0,2,0,2,6,9,8,9,10,12,12,11,12,12,13,14,14,12,12,11,11,11,12,11,10,9,8,8,8,5,0,0,0,1,0,2,8,9,8,9,7,6,7,7,7,8,9,10,11,10,7,4,2,2,1,3,3,8,8,7,8,6,0,0,0,0,0,3,9,8,8,4,2,1,0,0,1,3,6,8,8,7,4,2,1,1,1,1,2,4,7,7,7,6,0,0,0,0,0,2,9,8,6,5,4,4,3,1,2,3,4,6,8,6,4,1,3,7,7,5,5,4,2,4,4,2,0,0,2,1,0,0,8,8,5,1,5,10,19,12,8,3,5,7,8,8,2,7,10,13,11,7,5,6,7,1,5,8,1,1,2,12,2,0,6,1,4,6,6,7,7,8,8,7,2,1,7,0,9,8,6,6,6,7,5,5,7,2,8,8,2,2,5,19,2,6,8,2,8,7,5,3,3,3,2,3,8,1,5,0,8,6,4,5,4,4,6,8,6,4,9,9,2,2,4,19,3,4,7,3,8,10,7,4,5,7,6,7,8,1,17,4,5,7,5,6,5,7,9,8,8,4,9,9,3,2,3,19,13,4,5,7,7,9,8,6,7,7,7,9,8,4,17,14,6,7,10,8,8,9,10,7,10,9,9,9,7,4,6,19,19,7,4,10,10,6,8,10,9,8,9,9,6,8,17,15,3,6,7,8,8,8,8,8,11,9,8,9,7,5,6,19,19,14,7,10,5,8,8,9,10,10,9,8,1,11,17,16,8,2,9,9,9,9,9,14,9,8,8,9,8,7,18,19,19,18,7,10,9,8,8,7,9,9,9,2,7,13,19,18,10,7,3,6,13,14,5,8,8,8,8,8,8,19,19,19,19,19,19,11,9,8,4,13,11,7,5,3,12,11,14,13,10,11,3,4,5,5,5,7,8,7,8,2,14,19,19,19,18,19,19,16,9,8,6,5,5,5,6,4,6,4,6,5,2,3,6,7,6,5,6,8,8,7,8,2,19,19,17,19,18,19,19,18,9,8,7,6,6,7,10,9,3,2,1,1,2,7,9,12,11,8,8,8,8,8,8,11,15,19,19,19,19,19,19,19,9,8,8,7,7,10,10,8,8,7,5,6,8,7,7,9,10,9,8,8,8,8,8,17,19,16,19,19,19,19,19,19,12,9,8,8,8,8,7,6,9,6,7,7,4,5,6,6,7,8,8,8,8,7,8,18,17,17,16,19,16,19,19,19,19,8,9,8,8,8,6,4,2,2,3,2,1,1,1,4,6,7,8,7,7,7,9,19,19,18,18,19,17,19,19,19,19,8,7,8,8,7,5,5,5,7,9,10,8,6,8,7,8,7,7,6,6,6,16,19,15,17,19,19,19,19,19,19,18,18,6,6,7,7,8,8,7,5,4,4,5,7,7,8,7,6,6,5,5,8,17,19,19,15,19,19,19,19,19,18,19,17,12,5,5,6,7,7,6,4,3,3,3,5,6,6,6,6,6,5,4,11,19,18,19,19,18,19,19,19,19,19,19,19,19,12,5,5,6,6,5,5,6,7,7,7,7,7,7,7,6,4,5,14,19,19,18,17,16,19,19,18,18,19,19,19,19,14,4,5,7,7,7,9,8,7,6,8,8,8,8,6,4,3,6,14,18,19,16,19,14,19,19,16,19,18,18,19,19,15,4,3,5,8,7,6,7,5,4,5,5,6,4,3,2,4,7,15,19,18,17,16,19,17,19,19,19,19,19,19,4,2,6,4,3,3,4,3,3,3,3,2,3,2,2,2,3,6,7,12,19,19,19,19,16),(19,19,12,0,0,0,3,6,9,13,14,18,19,19,19,19,18,19,18,18,14,9,6,2,0,0,0,0,1,1,8,19,19,19,4,1,0,3,7,9,12,15,17,18,19,18,18,18,18,19,18,19,18,13,10,7,4,2,0,0,0,1,1,19,19,19,1,0,1,7,10,10,12,14,17,17,18,17,17,18,18,18,17,16,14,12,11,10,8,5,1,0,0,0,1,16,19,7,1,0,3,7,10,10,11,13,14,16,15,16,16,17,16,16,16,15,13,12,11,10,9,7,4,1,0,0,1,8,19,5,1,0,3,7,9,10,11,11,12,15,15,16,16,17,16,17,17,16,16,13,11,10,9,7,4,1,0,0,0,3,19,3,0,0,3,7,9,9,11,12,14,15,16,16,16,16,16,16,17,17,17,14,11,11,9,7,5,1,0,0,0,0,19,11,0,0,3,8,9,10,11,12,15,16,17,16,16,16,16,16,17,18,16,15,12,10,9,8,7,3,0,0,0,0,16,5,0,0,3,8,8,9,11,13,14,16,17,16,15,15,15,16,15,15,14,13,11,10,9,8,8,7,3,0,0,0,19,7,1,0,3,8,8,10,11,10,11,11,12,14,13,13,12,11,10,8,6,5,4,5,9,9,8,8,6,0,0,1,19,7,1,0,3,9,9,6,5,4,4,5,6,7,9,10,8,4,3,1,0,1,0,0,0,2,7,8,8,0,0,1,19,12,1,0,4,9,4,0,0,0,0,0,1,2,7,12,7,1,1,1,2,3,4,4,3,1,4,8,9,1,0,2,19,19,5,0,6,5,0,1,3,5,3,2,1,1,7,13,9,3,2,2,5,8,9,6,5,5,7,8,9,3,1,5,19,19,14,1,8,8,4,4,6,7,6,4,2,1,7,15,13,4,1,3,6,6,5,6,5,6,7,8,9,4,1,5,19,19,8,2,8,9,6,5,5,5,5,3,1,3,7,15,15,6,6,1,1,2,2,1,4,8,9,9,9,4,1,5,19,19,2,3,7,10,8,4,2,1,1,2,4,7,8,16,14,7,9,7,4,3,2,3,7,10,10,9,9,5,0,5,19,19,3,4,5,10,10,7,5,4,6,8,10,8,8,14,12,8,9,12,13,10,10,12,12,12,10,9,9,7,1,6,19,19,5,6,3,11,10,11,12,12,11,13,12,9,9,14,13,9,9,10,15,14,13,13,12,11,9,8,9,8,3,5,19,19,13,7,3,11,10,10,12,12,13,14,11,9,10,15,15,10,8,10,14,14,13,11,9,9,8,8,9,8,8,7,19,19,19,8,6,10,9,9,10,12,14,13,10,7,10,17,17,10,9,8,13,14,14,12,11,9,8,8,9,8,8,9,19,19,19,9,8,11,8,9,10,12,14,12,8,8,7,8,10,7,7,7,10,12,12,10,9,8,7,9,9,7,7,7,19,19,19,11,8,10,9,8,11,11,12,11,8,5,1,4,4,1,2,6,9,10,10,10,9,8,8,9,8,6,6,6,19,17,19,8,8,9,9,8,9,10,11,9,8,7,1,2,2,2,3,8,10,9,9,9,8,7,7,8,8,15,19,19,19,19,18,14,7,10,9,8,8,9,9,8,9,4,1,1,1,1,0,2,8,11,9,6,8,7,7,8,8,16,19,16,19,19,19,19,19,18,10,8,8,8,8,7,2,1,1,3,5,3,2,1,1,2,8,7,7,7,7,7,8,17,16,19,19,18,19,19,17,18,9,8,8,7,5,1,1,1,3,2,5,2,2,2,2,1,1,7,7,7,7,8,8,14,17,15,17,18,19,18,19,18,12,8,8,7,1,1,1,1,2,3,1,3,5,2,1,1,1,4,7,7,7,8,6,11,15,19,19,19,17,19,19,19,19,8,7,7,1,1,3,4,5,6,6,6,4,3,4,4,2,3,7,7,7,7,2,5,12,19,19,19,19,19,17,19,19,8,7,7,2,4,6,4,2,1,1,1,1,2,5,5,4,3,6,6,6,6,0,4,7,19,19,19,19,19,19,19,19,19,6,6,3,4,5,6,6,5,4,5,7,8,7,5,3,3,5,5,5,8,0,0,3,8,19,19,19,19,18,18,14,16,7,4,3,4,6,8,10,11,13,13,13,12,9,7,4,4,5,4,6,7,0,0,0,6,17,19,19,19,19,19,18,19,8,5,4,4,5,4,4,8,10,12,7,4,4,5,4,2,3,4,6,7,0,0,0,2,19,19,18,19,18,19,15,19,8,6,2,2,2,3,2,3,5,5,3,1,2,2,1,2,3,5,6,7,0,0,1,1),(19,3,1,1,1,0,0,0,1,1,0,1,1,2,3,3,4,5,6,7,5,4,4,3,2,0,0,1,1,1,3,19,5,0,0,1,0,0,0,0,0,0,1,2,4,5,6,7,9,10,10,10,9,8,7,6,4,0,0,0,1,1,1,2,0,0,0,1,0,0,0,0,0,0,2,4,6,7,9,11,12,13,13,14,12,9,8,7,5,1,0,0,1,2,1,1,1,0,0,0,0,0,0,0,0,0,4,7,8,10,11,12,13,13,13,14,12,11,9,7,6,3,0,1,1,1,1,1,0,0,0,0,0,0,0,0,1,3,7,11,13,14,14,14,14,15,14,14,12,10,8,8,6,3,0,1,1,1,1,1,0,0,0,0,0,0,1,4,5,8,13,15,15,16,15,15,15,15,15,15,13,10,9,8,6,3,1,1,1,1,1,1,0,0,0,0,0,4,6,9,11,14,17,17,17,16,16,15,16,16,16,16,14,12,9,7,6,3,1,1,1,0,1,0,0,0,0,0,2,6,8,11,12,14,14,15,15,15,15,15,15,14,14,12,12,12,10,9,7,5,1,0,0,0,0,0,0,0,0,1,5,7,8,8,8,8,8,9,9,12,12,11,11,10,8,7,6,5,5,4,6,6,3,0,0,0,0,0,0,0,0,2,6,6,3,3,2,2,1,2,5,7,8,8,7,5,2,1,0,1,2,3,3,4,4,0,0,0,0,0,0,0,0,4,6,4,3,3,4,3,2,1,1,3,6,7,5,2,2,2,4,7,7,5,3,3,4,0,0,0,0,1,0,0,0,5,5,4,5,7,11,12,8,3,3,3,7,12,7,3,3,5,9,12,10,6,5,4,4,1,0,0,0,0,0,0,0,5,5,4,4,5,9,10,8,4,3,4,10,19,13,5,3,4,7,9,7,5,4,4,5,2,0,0,0,0,0,0,0,6,6,5,4,5,5,5,4,2,3,7,10,18,16,6,3,2,3,4,4,4,3,5,6,5,0,0,1,0,1,0,0,7,6,6,4,1,1,1,2,4,7,8,12,17,17,8,7,3,2,1,1,2,5,6,7,6,1,0,1,1,2,0,1,7,7,8,7,5,4,5,6,9,12,9,11,15,17,10,8,9,5,5,4,6,6,8,8,7,3,0,1,2,8,1,1,7,7,9,10,9,9,9,9,13,13,8,11,17,19,15,8,12,11,9,9,9,10,10,8,7,4,1,3,16,19,2,1,7,8,10,11,13,13,13,14,15,11,7,11,16,19,15,10,9,13,13,12,12,10,9,8,7,6,4,7,19,19,8,2,7,8,9,10,12,15,15,15,13,9,10,9,11,13,10,8,10,11,13,13,12,10,9,8,7,6,5,18,19,19,19,6,7,7,8,10,12,13,14,14,12,8,6,2,3,4,2,1,5,10,11,11,10,9,8,7,6,6,8,19,19,19,19,10,7,7,8,9,10,11,12,12,13,10,3,2,3,2,2,2,4,9,9,9,9,8,7,7,6,7,10,19,19,19,19,16,7,7,8,8,10,10,11,12,12,9,8,7,6,4,6,6,6,8,9,8,8,7,6,6,5,6,8,19,19,19,19,12,8,6,7,7,8,9,10,10,9,9,9,9,10,12,10,8,7,7,7,7,8,7,6,5,5,6,8,19,19,19,19,16,6,6,6,7,8,8,8,7,9,8,4,3,3,3,3,3,4,7,6,5,7,6,5,4,5,9,19,19,19,19,19,19,19,7,5,6,7,8,7,5,3,1,3,4,3,2,2,1,1,1,4,5,7,5,5,5,5,19,19,19,19,19,19,19,19,8,5,5,6,7,6,4,5,6,7,12,12,10,11,8,5,4,3,4,6,5,4,5,6,19,19,19,19,19,19,19,19,18,5,5,5,5,4,5,6,5,3,3,3,3,3,3,3,4,4,4,4,4,4,4,12,19,19,19,19,19,19,19,19,14,5,4,4,4,4,4,4,3,2,1,1,1,1,1,2,3,4,3,3,3,3,4,19,19,19,19,19,19,19,19,19,19,19,4,3,3,3,4,3,3,3,3,3,3,3,2,2,2,2,2,2,2,3,19,19,19,19,19,19,19,19,19,19,19,19,12,3,2,2,3,5,4,4,4,4,3,3,3,3,2,2,2,1,2,5,19,19,19,19,19,19,19,19,19,19,19,19,19,19,2,1,2,3,3,3,3,2,1,2,2,3,2,2,1,1,2,5,16,19,19,19,19,19,19,19,19,19,19,19,19,13,3,1,1,2,2,1,1,1,1,1,1,1,1,1,1,2,3,6,0,19,19,19,19,19),(13,3,3,1,1,1,2,2,2,2,2,3,3,3,4,3,3,2,2,3,3,1,3,2,3,3,2,1,1,3,3,2,4,3,2,1,1,1,1,1,1,1,1,2,2,2,2,2,2,1,2,2,1,1,2,1,2,2,2,0,0,2,2,1,4,3,1,1,1,1,0,0,1,1,2,2,1,2,2,1,1,1,1,1,1,0,1,1,1,1,1,0,0,1,2,1,3,3,1,1,1,1,0,0,0,1,1,1,3,1,1,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,1,1,3,3,1,1,1,0,0,0,1,1,1,1,3,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,1,1,2,2,0,1,1,0,0,0,1,1,1,1,2,1,0,0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,2,2,1,2,1,0,1,0,1,1,2,3,1,0,1,0,0,0,0,0,1,1,0,0,0,0,2,0,0,0,0,0,1,2,1,2,1,1,1,1,1,1,1,2,2,1,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,1,2,0,1,0,1,2,2,2,2,3,4,5,5,5,5,5,4,3,3,3,4,4,4,4,3,5,2,0,0,0,0,1,1,1,0,0,4,8,7,6,5,4,3,5,6,7,9,9,6,5,4,4,5,6,8,6,7,7,6,0,0,0,0,1,1,1,0,1,6,8,8,7,6,5,5,5,5,9,13,11,7,5,3,4,6,8,10,8,8,8,7,5,3,1,0,1,1,1,1,4,7,8,9,10,10,7,4,3,4,11,19,19,11,3,2,3,5,6,8,8,7,8,10,9,7,1,0,1,0,0,2,7,8,7,7,7,6,5,4,2,5,12,19,19,12,6,6,2,1,1,1,2,11,11,11,11,9,4,0,0,0,0,3,10,11,9,5,6,4,1,2,6,9,12,19,19,13,13,10,8,11,9,10,11,12,13,13,11,10,5,0,0,0,0,5,12,14,14,10,8,8,10,11,14,15,14,19,19,13,13,15,18,10,12,15,14,16,15,13,11,9,4,0,0,0,0,5,13,16,15,16,16,15,12,15,15,14,14,19,19,15,12,14,18,19,18,17,18,19,15,13,9,9,3,0,0,0,0,4,13,16,18,19,19,18,19,19,15,14,14,19,19,15,13,13,17,19,18,17,15,14,12,10,9,8,3,0,1,0,0,3,11,13,15,17,17,19,19,18,15,12,15,19,19,14,12,10,14,18,18,16,15,13,10,9,8,6,2,0,1,0,0,1,10,12,12,15,18,18,18,17,11,14,13,15,15,12,12,10,9,16,15,14,13,11,10,8,7,5,2,0,1,0,0,0,8,11,12,14,16,18,17,14,10,11,8,8,7,6,7,7,9,9,13,13,12,9,8,7,7,4,3,0,1,1,1,0,6,11,11,12,15,15,15,12,11,6,1,4,5,3,2,6,13,13,9,11,10,9,7,7,7,3,3,0,2,2,1,0,4,9,10,11,13,14,13,15,14,4,3,4,3,3,4,13,14,15,12,8,8,7,6,6,6,4,3,0,1,1,1,2,3,8,10,11,12,13,14,14,13,13,10,7,5,8,11,12,12,12,13,10,6,6,5,5,5,4,3,1,2,1,1,1,2,6,8,9,9,10,11,11,12,13,12,11,10,11,11,10,9,9,9,10,8,8,7,6,6,4,2,0,1,1,0,0,1,6,7,7,8,10,9,9,8,10,11,12,17,9,8,9,8,5,5,7,10,9,7,6,5,4,1,0,2,1,0,0,0,4,7,8,9,7,6,6,8,6,3,2,3,3,4,3,2,4,2,6,10,10,7,6,6,1,0,1,2,0,1,0,0,3,9,9,11,10,6,3,5,6,8,11,12,11,10,10,10,10,9,6,9,9,7,7,5,0,0,1,3,1,1,0,0,1,7,10,10,11,10,11,10,10,9,6,5,6,7,8,10,11,10,10,8,7,7,8,6,4,12,19,7,6,1,1,0,0,8,10,10,9,10,11,10,10,9,9,12,16,17,15,12,11,10,10,9,8,8,7,7,15,19,19,19,19,19,2,1,1,7,9,9,9,10,11,12,12,13,19,19,19,19,18,14,12,11,10,10,8,9,8,6,5,9,18,19,19,19,19,19,19,19,9,10,9,10,11,12,13,16,16,18,17,17,15,14,12,11,10,8,7,7,6,4,5,0,1,19,19,19,19,19,19,19,18,8,10,9,10,11,12,13,13,14,13,13,11,10,10,9,7,6,6,6,4,4,4,0,0),(19,19,18,4,2,3,10,11,10,11,12,12,13,14,13,14,13,12,12,11,10,9,9,9,7,3,1,2,2,10,19,19,19,19,4,2,2,8,10,10,10,11,12,13,15,15,15,15,14,14,13,13,11,10,9,9,8,5,2,2,2,2,10,19,19,11,1,2,4,9,10,9,10,11,13,14,15,14,14,14,14,13,13,12,12,10,9,8,7,6,3,1,1,3,3,17,19,2,2,2,6,9,9,9,11,12,14,14,14,13,13,13,13,13,12,12,11,10,8,8,7,6,3,1,0,1,2,5,19,2,1,2,7,9,8,10,11,11,13,13,13,12,13,14,13,12,12,11,11,10,9,8,7,6,3,1,1,1,2,2,4,2,1,2,7,8,8,10,11,11,12,13,14,13,14,13,13,13,12,11,10,10,9,8,7,7,4,2,1,0,1,2,2,2,1,2,5,7,8,9,10,11,12,11,13,13,13,13,12,12,12,12,10,10,9,8,7,7,4,2,1,0,0,1,2,1,1,2,5,7,8,9,11,11,12,13,12,12,12,13,12,12,11,9,6,7,7,8,7,7,6,2,0,0,0,1,2,1,0,2,5,8,8,9,10,9,10,11,11,12,12,11,10,9,4,1,1,1,1,5,8,7,6,3,1,0,0,2,2,1,0,2,5,7,8,6,4,2,2,4,8,9,9,9,8,5,2,1,1,1,1,1,3,7,6,4,0,0,1,1,2,0,1,1,5,6,4,1,0,0,1,1,4,6,9,9,6,3,2,2,2,4,4,3,2,4,6,5,0,0,0,1,3,1,1,1,5,6,2,1,2,3,2,2,2,4,8,12,10,2,2,3,4,6,6,4,4,3,6,6,1,0,0,1,3,2,1,0,6,6,2,4,4,4,4,2,2,2,9,13,11,3,1,2,5,5,4,3,5,6,6,7,3,0,0,1,3,1,1,0,7,5,3,5,6,5,4,3,1,2,8,12,11,6,4,1,1,2,2,2,5,5,7,6,6,0,1,1,8,0,0,0,8,5,5,4,4,6,3,1,3,5,8,10,12,7,7,4,4,5,6,5,6,6,8,7,7,1,0,2,19,1,0,0,7,7,6,4,3,2,3,4,5,6,7,13,13,8,6,9,8,6,6,8,9,9,9,7,7,2,1,3,19,3,1,0,8,8,7,6,6,5,5,6,9,6,8,14,15,9,7,8,10,12,12,11,10,9,7,6,7,3,1,2,19,13,1,0,7,8,8,7,8,8,9,11,9,7,9,14,13,10,7,6,10,11,11,10,9,7,6,6,6,5,2,4,19,18,8,1,5,8,8,9,10,10,12,11,8,7,8,14,11,8,6,6,6,8,10,9,8,6,6,5,6,6,5,5,19,19,17,1,2,8,8,9,9,10,12,10,6,6,6,7,7,5,2,4,4,6,7,7,7,6,5,5,6,6,5,7,19,19,18,5,4,8,7,8,9,9,10,8,6,4,2,3,3,2,1,3,6,7,5,6,6,6,5,5,6,6,6,7,19,19,19,8,4,8,7,7,8,8,8,7,7,7,2,2,1,2,4,5,5,7,7,6,6,6,5,6,6,6,7,7,19,18,18,12,7,8,7,6,7,7,7,6,6,6,5,4,2,4,5,6,5,5,7,6,6,5,5,5,5,6,4,6,18,19,19,16,8,8,7,6,6,7,6,7,6,5,6,5,4,4,5,5,5,5,5,5,6,5,5,5,5,6,12,12,19,19,19,16,8,8,7,6,6,6,4,6,5,5,6,7,8,8,5,3,3,5,4,5,5,5,5,5,5,6,13,13,19,19,18,19,18,8,7,6,6,5,6,5,5,5,3,1,1,1,0,0,2,1,1,3,5,5,5,5,5,5,12,15,19,18,19,16,19,19,7,6,6,7,5,2,2,2,4,5,6,6,7,7,5,4,4,5,5,5,4,5,5,6,16,14,19,19,19,16,18,19,8,7,6,6,5,5,5,5,6,7,6,5,4,3,3,4,6,5,5,4,4,4,5,14,13,13,19,19,19,19,19,19,10,7,6,5,5,5,7,5,3,3,2,2,2,3,5,6,5,5,4,4,4,4,4,14,15,14,19,19,19,19,19,19,17,6,6,5,5,6,6,6,6,5,4,4,5,6,7,6,5,5,4,4,4,4,4,5,12,16,19,18,18,19,19,19,19,7,5,5,5,5,5,7,8,9,10,9,8,9,8,6,5,5,4,4,4,3,5,0,13,16,19,19,19,19,18,19,18,4,5,5,5,5,6,7,7,7,8,7,7,7,6,5,5,4,4,3,2,4,5,0,1,14),(0,1,1,0,0,0,0,0,1,1,3,4,5,6,5,5,4,3,5,5,3,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,1,1,3,5,7,8,9,8,8,8,7,9,8,8,7,4,2,1,0,0,0,0,0,0,0,0,1,0,1,0,0,1,3,4,6,7,8,10,9,9,9,10,10,10,9,9,8,7,6,3,2,1,1,0,0,0,0,0,1,0,1,0,0,2,4,6,7,8,8,10,10,10,10,11,12,11,10,10,10,9,7,6,4,3,1,0,0,0,0,0,1,1,0,0,0,2,6,7,7,8,9,11,12,11,11,11,12,11,10,11,11,9,7,6,5,4,2,0,0,0,0,0,1,1,0,0,0,4,6,6,6,7,9,11,13,12,12,12,12,12,11,12,10,9,7,6,5,4,2,1,0,0,0,0,1,1,1,0,2,5,6,7,8,8,10,11,12,13,13,13,13,13,13,12,11,9,8,7,5,5,4,2,0,0,0,0,1,1,0,2,6,6,7,7,8,9,9,10,12,12,12,13,12,11,11,11,11,9,8,8,7,6,5,4,4,0,0,0,1,1,0,6,6,6,4,2,2,2,2,4,5,7,9,9,10,10,7,6,6,5,4,3,2,3,5,5,5,0,0,0,1,1,0,7,6,4,5,4,5,3,3,6,6,4,6,7,7,6,5,4,5,5,2,2,2,2,2,5,5,1,0,0,2,1,1,7,6,9,6,4,4,3,2,3,3,3,2,5,5,3,1,2,2,2,3,4,3,4,4,4,5,1,0,0,5,2,3,5,5,10,8,10,9,10,9,6,4,3,5,10,7,6,4,6,3,4,7,7,7,6,6,6,4,0,0,2,5,7,9,7,6,11,6,6,6,6,5,3,3,4,3,4,5,3,3,3,2,7,7,5,6,8,5,5,3,6,4,4,8,7,6,6,7,7,6,4,2,2,2,2,3,4,2,11,12,4,4,2,2,2,3,2,3,5,6,6,6,6,5,4,9,6,5,5,5,7,8,7,3,3,2,4,5,8,5,14,15,8,3,5,4,3,2,3,4,6,7,6,4,4,4,6,5,2,4,5,7,7,10,9,6,6,6,6,5,3,8,14,16,9,3,5,7,6,5,6,8,11,7,6,4,5,2,5,5,7,11,8,11,8,8,6,6,6,7,5,5,5,8,15,17,9,7,2,7,8,7,7,7,7,7,6,7,8,7,4,8,7,6,8,7,14,7,8,8,8,8,5,3,8,11,16,18,10,8,3,4,7,7,7,7,6,7,9,5,6,9,7,6,10,7,8,8,7,5,4,4,4,4,3,8,14,12,17,19,11,12,12,4,3,9,7,7,7,12,6,7,5,9,5,12,7,6,8,8,7,4,4,4,5,7,8,10,11,10,13,13,9,9,9,6,5,3,3,3,3,4,6,7,5,5,8,19,11,8,10,8,6,5,5,7,7,8,8,6,2,3,6,6,3,2,4,6,7,5,3,3,3,4,6,7,7,8,19,19,17,11,7,8,6,5,5,5,6,7,6,5,1,2,2,2,1,0,3,5,5,4,4,3,3,4,6,5,8,10,19,19,19,18,19,8,6,5,5,5,5,5,4,3,1,1,0,0,0,0,1,2,2,3,4,3,3,4,6,19,13,19,19,19,19,19,19,8,6,5,5,4,4,3,1,1,0,0,0,0,0,0,0,1,0,2,3,4,4,5,6,19,19,19,19,19,19,19,19,9,6,5,5,4,3,2,0,1,1,2,2,2,2,2,2,1,0,1,3,4,4,5,7,19,19,19,19,19,19,19,19,16,7,5,5,3,2,1,1,1,2,3,3,3,4,3,2,1,0,1,2,4,4,5,13,19,19,19,19,19,19,19,19,19,6,6,5,3,2,2,3,4,5,5,5,5,5,6,4,3,2,2,2,4,4,5,18,19,19,19,19,19,19,19,19,19,13,5,5,4,3,3,3,4,4,4,4,3,3,4,4,3,3,3,3,4,4,6,19,19,19,19,19,19,19,19,19,19,19,6,5,4,4,3,3,4,3,3,2,2,2,3,3,3,3,4,4,4,4,6,19,19,19,19,19,19,19,19,19,19,19,8,5,4,4,4,4,5,5,5,4,4,4,4,4,4,3,3,4,4,3,6,19,19,19,19,19,19,19,19,19,19,19,9,4,4,4,4,4,5,5,7,7,7,6,5,5,4,4,4,4,3,4,6,19,19,19,19,19,19,19,19,19,19,19,9,5,2,4,5,4,4,4,5,5,5,4,4,4,3,4,4,3,3,4,6,19,19,19,19,19),(19,4,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,3,2,3,3,3,1,0,0,0,0,1,0,1,1,19,1,0,0,0,0,0,0,0,0,0,1,1,2,3,4,5,6,4,5,6,6,4,3,2,1,1,1,0,0,0,0,11,0,0,0,0,0,0,0,0,0,1,2,4,5,7,8,8,7,8,8,8,7,5,4,3,2,1,1,0,0,0,0,1,0,0,0,0,0,1,0,1,2,3,4,6,8,10,10,10,9,9,10,9,7,6,5,5,3,2,2,0,0,0,0,0,0,0,0,0,0,1,2,4,4,4,5,9,10,11,11,10,11,11,11,9,8,7,6,5,4,3,2,1,0,0,0,0,0,0,0,0,2,2,5,5,5,6,8,11,12,11,13,12,12,12,11,10,9,7,7,6,5,4,2,2,0,0,0,0,0,0,0,1,2,4,5,5,6,8,10,11,12,13,13,13,13,12,11,11,10,9,7,7,6,5,3,3,0,0,0,0,0,0,0,2,3,5,6,7,8,10,11,11,11,13,13,13,13,10,11,11,11,11,9,6,6,5,4,3,1,0,0,0,0,0,0,4,5,6,4,4,5,5,5,6,9,9,11,11,10,9,8,5,4,4,4,4,4,5,5,4,2,0,0,0,0,0,0,5,5,4,4,4,4,4,4,4,4,7,9,10,8,5,4,4,5,6,7,6,4,4,5,5,4,0,0,0,0,0,1,5,5,5,7,8,11,10,8,5,5,6,9,8,7,6,5,7,10,11,12,9,7,5,6,6,5,1,0,0,0,0,2,6,6,6,7,8,11,11,9,7,6,7,10,10,8,6,7,8,9,10,12,9,7,6,6,6,5,1,0,2,0,0,3,7,6,7,6,7,8,8,6,6,6,8,12,13,9,7,5,6,8,9,9,7,6,6,6,7,6,2,0,5,0,0,4,8,6,3,2,1,1,1,2,4,8,8,12,14,8,7,6,3,1,2,3,3,4,4,6,6,6,2,0,11,0,0,6,8,8,8,6,4,3,3,6,8,10,10,12,14,7,9,8,6,3,3,3,3,4,6,7,8,7,1,0,15,6,1,7,8,9,9,11,12,12,11,11,12,11,10,13,14,8,9,11,11,10,11,10,10,9,9,8,8,8,1,0,7,2,4,8,8,9,11,12,14,13,13,13,12,10,10,13,13,10,9,12,14,14,14,14,14,13,11,10,8,8,1,3,12,4,4,8,8,9,11,13,14,14,14,15,11,9,10,12,11,10,10,11,13,15,14,14,14,14,11,9,8,8,2,5,19,7,6,8,7,8,10,11,12,14,14,12,8,9,10,12,11,10,8,8,12,14,15,13,13,12,10,8,7,8,3,4,19,10,4,8,6,7,9,10,11,12,12,8,10,11,9,10,10,9,11,8,9,12,13,12,12,11,9,7,7,7,5,4,19,13,5,9,6,6,8,8,9,10,8,7,7,5,4,4,4,4,7,6,7,9,10,10,10,9,8,7,6,7,8,4,18,16,8,8,6,6,6,7,7,7,7,7,3,2,2,2,2,2,2,3,7,7,9,8,8,7,7,6,6,7,7,7,19,19,10,9,6,6,6,6,6,7,7,7,7,5,5,5,4,4,4,6,7,7,7,7,7,7,6,5,6,7,8,7,18,19,16,8,7,6,5,5,6,6,6,6,6,7,8,9,9,9,8,8,8,7,7,6,6,6,5,6,6,7,8,12,19,19,19,16,8,6,5,5,5,6,5,5,7,8,7,9,8,7,9,7,6,6,5,5,5,5,5,5,6,7,10,18,19,19,19,19,13,6,6,5,5,5,4,3,3,3,3,3,3,3,3,3,3,5,5,5,5,5,5,5,6,11,19,19,19,19,19,19,19,7,6,5,6,5,3,4,4,6,9,8,8,8,6,5,4,4,6,6,5,5,5,5,6,15,19,18,19,19,19,19,19,8,6,6,6,6,7,7,6,5,4,4,4,4,5,6,7,7,6,6,6,5,5,5,7,17,19,19,19,19,19,19,19,9,7,6,5,5,6,7,6,6,5,4,5,6,6,7,6,6,5,5,4,4,4,5,8,19,19,18,19,19,19,19,19,17,7,6,5,5,6,7,7,8,9,10,10,9,8,7,6,6,5,4,4,4,4,5,17,19,19,19,19,19,19,19,19,19,7,6,5,6,6,6,7,8,10,10,10,9,8,7,6,6,5,4,4,4,5,9,19,19,19,18,19,19,19,19,19,19,7,6,6,6,6,6,7,8,9,8,9,9,8,7,7,5,5,4,4,5,5,15,19,19,19,19),(9,1,0,0,0,0,3,7,10,10,10,7,3,2,3,4,7,13,15,16,15,14,12,11,9,2,0,1,0,0,2,19,19,1,0,0,0,4,9,11,11,12,13,12,11,10,10,11,15,16,17,17,15,14,12,11,10,6,1,0,0,0,2,19,19,0,0,0,2,9,11,11,12,13,15,16,16,15,15,15,15,15,16,17,15,14,12,11,10,8,3,0,0,0,2,19,19,0,0,0,6,9,10,12,12,13,14,16,15,15,15,14,14,15,15,15,15,13,12,11,10,8,5,0,0,0,3,19,19,1,0,0,7,10,10,12,12,13,15,16,16,16,16,16,15,16,16,15,15,13,11,11,9,9,6,1,0,0,1,19,19,2,0,0,6,9,9,12,12,14,15,17,17,17,17,16,16,17,17,16,15,13,12,11,9,8,7,1,0,0,2,19,19,2,0,0,5,9,9,11,12,14,16,18,19,18,16,17,17,17,18,18,15,14,13,11,9,8,7,0,0,0,4,19,19,2,0,0,4,9,9,11,13,13,15,16,16,17,18,17,17,17,16,16,14,13,12,11,10,8,8,0,0,0,8,19,19,3,0,0,7,9,10,10,10,10,11,12,12,13,15,16,13,12,12,12,11,9,7,7,9,9,8,1,0,0,12,19,19,7,1,0,9,9,5,2,3,2,2,4,5,6,8,10,9,7,5,3,2,1,1,1,1,5,8,4,0,0,11,16,19,7,1,1,10,4,1,1,2,1,1,0,0,1,4,5,5,3,1,0,0,1,2,2,2,1,6,8,0,1,7,19,18,5,2,3,10,5,4,4,5,6,4,3,2,2,4,6,7,4,2,2,3,5,5,4,4,4,7,9,1,4,3,13,16,6,2,7,11,7,5,4,6,7,7,4,2,2,5,16,18,7,1,1,3,7,7,6,6,6,7,9,1,5,5,10,16,8,8,12,11,9,7,5,2,2,1,0,2,4,10,16,18,9,4,2,0,1,1,1,5,7,9,10,6,8,8,12,19,11,8,12,11,12,10,9,6,4,4,4,5,11,11,13,18,9,10,5,3,4,4,6,9,11,10,10,9,6,9,14,18,11,6,12,12,11,12,12,10,8,8,9,12,11,9,14,19,9,10,11,9,8,9,11,11,12,10,10,9,6,9,18,19,11,8,11,12,12,14,15,15,16,15,16,12,11,10,13,19,10,9,10,14,15,13,14,13,12,10,10,8,8,10,13,19,11,11,10,11,11,13,15,17,17,18,16,12,7,10,13,19,11,8,9,14,16,16,14,12,11,10,8,8,10,8,19,19,14,10,10,9,10,12,15,17,16,16,15,10,10,11,13,17,11,10,6,12,14,15,14,11,9,9,9,7,8,10,16,19,19,12,12,9,10,11,12,14,17,15,14,8,9,11,13,14,12,9,7,9,12,14,13,11,9,7,7,9,10,11,19,19,19,8,6,8,9,10,10,12,13,13,10,8,5,3,6,8,6,3,6,6,9,11,11,10,8,6,7,6,7,16,19,19,19,18,19,9,9,9,10,10,10,10,7,8,8,3,4,3,2,3,8,7,8,8,9,9,8,7,7,16,15,19,16,19,19,18,19,12,9,8,9,9,10,8,9,9,8,7,4,3,5,7,8,8,8,8,8,7,7,6,7,18,19,18,19,18,19,17,19,18,9,8,8,8,8,8,8,8,9,10,9,9,10,10,7,7,7,8,7,7,6,6,8,17,19,19,18,19,19,19,16,19,8,8,7,8,8,6,3,4,2,2,3,3,2,1,2,2,5,8,8,7,6,7,16,15,19,15,19,19,18,19,19,19,8,7,7,7,8,5,5,6,4,5,2,1,4,6,5,6,4,7,7,7,6,7,19,19,19,18,16,18,19,19,19,19,17,7,7,7,6,6,7,7,5,6,8,8,6,4,4,7,5,5,6,7,6,10,19,19,19,16,18,19,19,19,19,17,19,5,6,6,6,6,6,7,5,3,2,2,2,3,6,7,5,6,6,6,5,14,19,19,18,19,17,19,19,17,19,19,10,6,4,5,5,6,6,6,6,3,2,2,2,4,6,6,6,6,5,4,6,2,14,14,17,19,19,18,19,17,19,15,2,8,4,3,4,6,8,9,9,10,12,12,11,10,9,8,7,5,4,3,7,1,5,18,17,18,16,19,19,19,19,11,1,8,6,3,3,4,7,9,10,12,12,9,11,11,9,8,6,3,2,4,8,0,3,18,18,16,17,19,19,19,19,5,1,8,6,4,3,3,3,7,8,8,6,3,6,6,6,5,2,2,3,5,8,0,2,10,15,19,19),(8,7,6,6,5,5,6,7,9,11,9,9,9,10,7,8,9,6,6,7,6,6,5,5,5,5,4,4,5,4,5,5,6,5,5,5,5,4,4,8,12,13,13,12,10,10,10,6,8,7,8,6,7,7,4,4,4,5,5,6,6,4,3,4,4,2,3,4,4,4,6,12,13,13,12,14,11,10,10,8,8,8,8,8,7,6,5,6,6,7,5,4,4,4,4,4,4,2,1,2,4,6,9,12,13,14,14,12,12,8,8,8,8,10,9,8,7,8,6,5,5,7,5,3,3,3,3,4,5,2,2,3,4,7,11,12,13,14,13,13,12,9,9,7,7,10,12,11,9,7,6,5,5,5,4,3,1,2,3,3,3,2,2,3,4,6,10,13,14,14,14,14,12,12,7,8,8,9,10,10,11,8,7,6,5,4,3,3,3,1,2,3,3,2,2,2,3,5,10,13,14,15,15,15,15,12,9,8,9,11,11,12,12,11,9,8,7,5,2,2,1,3,2,3,4,2,1,1,2,5,11,14,15,16,15,15,14,14,11,8,9,11,13,15,12,11,10,9,7,6,2,1,1,1,2,2,1,1,0,2,3,6,13,16,17,16,15,14,13,13,12,10,8,11,13,13,12,12,12,10,10,7,2,1,1,1,3,0,2,0,1,3,1,9,13,15,14,13,11,9,11,10,11,10,10,11,12,12,13,14,15,13,11,8,4,0,1,1,2,1,2,2,2,2,1,11,12,9,7,4,3,3,4,6,7,8,10,9,7,6,6,5,7,9,10,9,5,0,1,1,1,2,3,2,3,0,3,12,8,6,5,7,6,3,2,3,5,13,13,6,3,2,1,2,3,4,5,9,6,0,1,0,1,3,6,3,3,0,9,12,9,6,7,8,8,4,2,2,5,19,19,7,2,1,2,5,4,4,3,5,8,2,0,0,1,2,13,7,4,1,11,13,12,9,5,5,4,5,6,7,11,19,18,10,5,3,2,2,3,5,4,6,8,5,0,0,0,3,19,17,5,2,13,14,14,14,12,11,12,13,12,15,12,19,18,10,13,9,7,7,6,6,8,9,10,8,0,0,1,3,19,19,7,5,13,15,17,18,18,19,19,19,18,15,12,19,16,10,13,16,17,16,14,13,13,13,12,9,1,1,2,3,19,19,8,8,12,14,17,19,19,19,19,19,17,14,14,18,16,11,12,15,19,19,19,18,17,14,13,10,3,2,3,6,19,19,8,10,12,12,15,16,19,19,19,19,13,11,14,19,19,12,10,13,19,19,19,18,16,14,12,10,7,2,7,19,19,19,11,10,12,12,14,15,18,19,19,18,10,14,13,16,15,12,13,10,17,19,19,17,14,12,10,10,9,1,17,18,19,19,11,12,12,12,13,14,15,17,17,15,9,7,6,8,6,5,9,9,15,16,16,14,12,11,10,9,9,2,18,19,19,19,12,13,11,12,12,12,13,14,14,15,12,2,1,3,2,0,1,11,14,13,13,12,11,10,10,9,9,6,16,19,19,19,19,13,11,11,11,11,13,14,16,13,10,10,8,3,3,8,8,10,13,13,12,10,9,9,9,9,9,7,19,19,19,19,19,8,11,10,11,11,14,14,15,12,11,12,10,8,7,11,10,10,11,13,12,10,10,9,9,9,9,14,16,19,19,19,19,3,11,10,10,11,14,13,12,11,11,8,10,15,15,9,10,10,9,11,12,11,10,8,8,9,5,19,19,17,19,19,19,16,11,10,10,12,14,14,6,4,3,2,3,2,2,3,4,4,5,8,11,12,10,8,8,8,17,16,19,19,19,19,19,18,15,10,10,12,14,12,9,9,7,9,10,10,8,8,7,4,3,5,9,11,10,8,8,8,19,19,18,19,19,19,19,19,19,10,10,11,12,11,12,13,12,10,6,5,4,6,8,10,11,11,9,10,9,8,8,9,19,19,19,19,19,19,19,19,18,9,10,10,10,11,10,11,10,8,7,6,5,7,8,9,10,10,9,8,8,8,7,19,19,19,19,19,19,19,19,19,19,12,9,10,9,9,11,10,9,9,7,6,6,7,8,8,8,8,9,8,8,8,7,19,19,19,18,19,19,19,19,19,19,14,9,9,9,10,12,13,14,17,18,18,17,16,12,10,10,9,8,8,8,7,19,19,19,19,19,19,19,19,19,19,19,14,10,7,8,8,12,14,15,18,18,14,16,19,16,15,12,9,7,7,6,17,19,19,18,19,19,19,19,19,19,19,19,14,11,7,6,7,9,11,12,12,12,11,12,13,12,12,10,8,6,5,6,18,19,19,19,19,19,19));
			yp_2D := ((358618,32481,-34093,-1293,-12380,6524,-286,3565,7133,2530,-10668,4403,-8857,615,5075,-6207),(358618,32481,-34093,-1293,-12380,6524,-286,3565,7133,2530,-10668,4403,-8857,615,5075,-6207),(362554,14827,-40549,5547,-8698,4842,1503,-3603,-2147,3467,-24138,11038,2122,3889,-8675,-10382),(242711,112871,1011,-35792,-13533,-26272,-14294,15053,-4706,7280,-17352,8090,-16496,-3951,-1821,-20862),(368447,33352,-68347,10329,-8691,13234,4388,-9447,764,2820,-23729,17678,-7885,-1670,-10763,-17588),(362555,51294,-63569,5558,-14105,17527,279,3805,9029,-16283,-12220,-7556,-25573,-8453,10007,-13853),(189641,-75444,-72649,46257,-195,53639,25845,10942,18327,-13186,-11121,-3398,-14398,-5229,-2531,-4349),(359405,18631,-59993,12182,-3080,17480,5032,-7701,2537,-3897,-15486,9985,-21992,-6339,-7368,-22083),(368746,35387,-31957,-3846,-19767,10758,7660,-15489,902,4643,4977,12819,269,9576,-1275,7236),(363140,49529,-29702,-7949,-26172,2959,3474,1480,4344,3909,-646,312,5009,4248,2914,8477),(369926,-21363,-7559,2700,3833,14391,10992,7260,-12136,3679,-42388,12684,-7970,-2460,-12944,-12815),(285041,8036,46385,-23170,-7729,-4950,5036,9625,1009,-4598,4662,-14939,-3748,1283,7382,7038),(294921,-746,48540,-23294,-10288,-4595,11710,-2199,-2735,7083,1795,6449,16054,3526,-4842,13856),(276021,102180,45189,-50173,-9841,-38957,-17260,12629,-15617,12045,-25545,5408,-6556,-5349,-8641,-10950),(288233,-6557,33914,-13327,3933,-9836,-3338,16823,-4644,-5915,-10519,-16760,-17132,-9363,4311,-6345),(288233,-6557,33914,-13327,3933,-9836,-3338,16823,-4644,-5915,-10519,-16760,-17132,-9363,4311,-6345),(270554,-92181,-25567,31674,6869,32512,23550,1213,1753,-401,-20090,7090,-503,-2387,-9082,-3355),(292660,7580,40470,-20748,-4819,-8502,-104,7488,-650,-5190,-407,-15755,-4660,-85,6691,6581),(290925,-14447,36335,-16745,-11826,9059,27470,-45645,-18187,13632,16690,34215,32818,6292,-21740,21984),(298664,24511,59040,-33779,-17500,-1984,10088,11771,5081,-2593,12290,-11227,5371,4853,6783,17755),(253354,31778,-72,-11671,-1403,-36493,-32848,23745,-2360,8931,-10686,-13967,6434,10244,10482,-3254),(293687,-22519,49586,-17862,9572,-28637,-23284,25269,-5244,24027,-30456,514,19737,24549,-1030,1097),(318827,4707,5092,-5471,8221,-34841,-39188,30926,-4780,-1958,-19601,-28836,-8204,7655,14519,-13390),(204643,91504,28865,-39206,-5103,-49938,-33085,18990,-11638,13459,-18459,-3171,-3773,1503,3785,-14994),(334520,1713,-3935,-1748,9916,-34048,-38179,21449,-9135,1924,-21217,-24243,-6062,4072,8280,-12891),(334520,1713,-3935,-1748,9916,-34048,-38179,21449,-9135,1924,-21217,-24243,-6062,4072,8280,-12891),(145765,-66968,-56936,38942,4681,28542,5481,17499,12434,-5805,-11144,-11032,-6128,7763,1238,-4265),(319713,15455,-10131,-2494,5224,-28543,-37475,25291,-3637,-6404,-14446,-33485,-14413,873,16304,-14365),(315022,-2221,-29761,7843,238,-35678,-30788,-16876,-14512,20318,3598,4978,20248,7123,-4818,9165),(317457,28584,16495,-17592,-673,-33724,-35396,33397,-5133,6573,-21740,-24755,-3405,13514,12782,-4354),(273219,-21849,-39478,16987,9730,-20040,-11605,471,-11458,19989,-10707,22342,3804,-36,-22788,-24859),(260141,-39930,-11147,9398,298,-16133,4045,-29190,-13097,34400,8989,45906,35607,2515,-27268,8735),(255264,-48717,-37966,22940,10323,-15068,-6198,-21242,-18120,28244,-8851,37805,18821,6225,-24871,-5683),(260742,111512,-5544,-34847,-22472,-47815,-23066,-2538,-9663,26652,-2593,19978,25558,8420,-12894,3131),(266266,-33222,-33581,16895,3688,-28763,-14628,-20760,-11038,33240,8226,32825,32166,4829,-20171,3776),(252581,-43362,-38610,21050,6156,-23706,-8876,-24850,-12475,37588,-2904,43069,35271,10437,-27184,4353),(157624,-85573,-63810,45933,5791,22813,8196,8386,11767,6773,-10395,3805,7377,6875,-8631,-52),(252581,-43362,-38610,21050,6156,-23706,-8876,-24850,-12475,37588,-2904,43069,35271,10437,-27184,4353),(257938,-24914,-28400,10275,-9539,-16147,5181,-42153,-12112,41187,14854,56826,57788,16946,-29673,25077),(240342,-39368,-36359,20329,9962,-32403,-18629,-11127,-17222,36425,-4401,32067,25514,5636,-24332,-7887),(268055,16483,31323,-21920,-20548,28167,46333,-39787,-2217,-2703,32765,38428,2540,4250,-14577,1661),(277085,-20504,41332,-13814,-6280,73885,75519,-35804,838,-35797,16183,22695,-44617,-15858,-16153,-21874),(308675,2409,60235,-27861,-17455,53380,59965,-23651,6180,-30851,26843,11399,-28654,-15001,1684,-1182),(265926,120786,57157,-62013,-28972,-5983,22225,-13427,-5016,10981,8011,33301,-69,2629,-16128,1184),(310832,5680,53265,-27127,-21131,72307,81095,-43930,4204,-31533,35880,30269,-29680,-11919,-8961,-4530),(296637,-4204,43847,-19472,-12236,70305,70662,-31300,4073,-36522,22895,17760,-45857,-16269,-8990,-14651),(154412,-71117,-38538,32729,-4202,60909,41465,4800,17970,-19148,2782,-2174,-17788,-2707,352,2392),(300185,11992,56537,-29096,-18269,52964,55462,-17593,8752,-28944,27058,8794,-33215,-14148,5421,563),(292649,-15030,39118,-14371,-7737,59621,62258,-27606,1718,-31685,18687,16342,-40396,-14394,-12111,-14490),(285020,-1097,40860,-18673,-12428,56631,57866,-21982,6419,-31110,23563,8818,-42109,-15581,-2381,-9709),(365383,8019,-69966,20610,-9334,24335,-4005,39959,20274,-22604,-24257,-31808,-27168,-2555,18115,-12601),(226446,-8068,-16786,8345,1738,6872,-7922,30003,10878,-24111,-3693,-32006,-32773,-13245,19738,-12129),(244500,-2610,-21010,8338,-479,10672,-6314,30284,12531,-29832,-6879,-34898,-35286,-14745,21435,-10411),(326646,120193,-4886,-36443,-15095,-30775,-28626,35316,-679,-832,-33361,-11274,-14849,61,7704,-11456),(248584,-7907,-21649,9653,1372,654,-13843,21211,8573,-20885,-2882,-28387,-24496,-10222,19185,-7329),(248584,-7907,-21649,9653,1372,654,-13843,21211,8573,-20885,-2882,-28387,-24496,-10222,19185,-7329),(266399,-88188,-55861,43716,694,25538,6459,33109,21173,-5556,-9289,-31020,-1377,6720,14104,6234),(241403,-10788,-12142,6645,1768,-9987,-19019,20582,6836,-12173,-327,-29271,-11883,-7122,17883,620),(231997,-4684,-14679,6451,2542,7390,-8461,22407,8217,-28087,-393,-32286,-35696,-15316,22289,-9021),(219627,-7994,-22628,10310,-289,-10472,-16243,15852,2545,-10501,4622,-20011,-14376,-10591,10920,-3404),(198159,-13347,10392,-277,6730,-33456,-21616,1614,-12227,-2183,23386,-11287,-5278,-10221,9178,-7688),(254176,-72507,25665,9845,23463,12071,11629,-11402,-12242,-26301,11641,-895,-38433,-32222,-2373,-34166),(272805,-63529,24031,8060,21992,-18572,-12738,355,-14838,-13264,7365,-9292,-20319,-25073,729,-24854),(135895,43215,26603,-22193,3449,-36709,-20567,9125,-13323,542,9213,-4969,-18243,-15981,3590,-23643),(267631,-36624,39825,-5592,10849,-31143,-19003,12156,-7875,-7504,24425,-19323,-8023,-15548,14192,-6604),(267631,-36624,39825,-5592,10849,-31143,-19003,12156,-7875,-7504,24425,-19323,-8023,-15548,14192,-6604),(119927,-58162,-12928,21815,4720,10735,2058,16458,9380,-14715,15637,-19783,-11098,-6543,13175,-530),(248616,-46963,17856,7208,19055,-7167,-10947,16612,-4168,-24245,22918,-25637,-43065,-28497,15818,-31923),(244184,-87557,-20287,28809,21190,10335,13774,-37594,-30454,4934,6817,34879,-5738,-11362,-21230,-23486),(259674,5494,57230,-24881,-7066,-17361,-6016,15968,431,-13309,28789,-24587,-4557,-10049,22689,9306),(335189,-44341,-12922,11318,2647,-4799,-2099,15538,1336,23085,-26407,19385,16508,12367,-9682,741),(315809,-35720,44872,-11294,9825,-5313,-9607,50150,8487,6149,-30328,-13715,-11870,12844,8,-13076),(326657,-11777,42930,-19705,-16410,-230,16270,-914,8135,19234,3434,22472,26844,6646,-15632,22926),(291787,62112,41372,-39306,-7346,-45352,-21813,16498,-14224,43015,-23417,21848,14750,15749,-20890,271),(326378,-32294,19044,-4070,-21,-17871,-7842,15654,-2216,27026,-13268,19175,19848,6508,-12415,10600),(315809,-35720,44872,-11294,9825,-5313,-9607,50150,8487,6149,-30328,-13715,-11870,12844,8,-13076),(250624,-73687,3927,13269,-8333,3698,8177,21032,11497,36925,-2583,17522,41123,27499,-7797,31572),(325312,6110,45627,-25070,-20384,7534,21994,-3215,13628,8562,18538,10132,16722,4212,-6290,24290),(295567,-25619,16240,-5584,-5301,-15536,3815,-17140,-7193,29801,-4491,38409,35545,12012,-22707,18297),(314133,-28552,20585,-7538,-10654,-13105,10168,-13172,-3901,39948,-790,44058,42347,11613,-30099,20233),(361462,-27801,3565,329,2365,45405,31128,-21533,-10128,-23104,-28409,16397,-18406,-4948,-7844,-10046),(323827,-20948,57734,-21094,1717,31991,25576,-10717,-1746,-25841,-11994,-3723,-14928,-5003,5938,-10),(327963,262,57794,-28533,-13227,44493,39962,-29902,-641,-32440,4083,4045,3640,1605,6686,12810),(268577,127026,65458,-66729,-20374,-28658,-3528,-9764,-16943,11116,-11299,20687,7982,2133,-10798,5130),(325850,21361,56543,-34010,-16465,42199,33267,-19345,5565,-32697,2685,-9890,-1177,4614,15177,21319),(325850,21361,56543,-34010,-16465,42199,33267,-19345,5565,-32697,2685,-9890,-1177,4614,15177,21319),(233624,-80505,-37727,33298,-4719,59736,33484,13217,21700,-20938,-14927,-14143,-3924,2895,5479,10596),(294696,12168,50748,-26454,-1370,10964,2950,29473,8414,-23366,-23082,-29119,-18096,-807,22891,-1813),(329420,-23673,42434,-15655,-1102,58155,45675,-40724,-8135,-32717,-3656,13895,-19401,2927,5039,153),(323404,44480,49817,-38300,-32566,28553,30220,-7862,16677,-10068,18701,-6018,13651,5224,6888,33734),(273948,26463,-14173,-3515,2584,-22146,-22329,20330,-741,-8639,-1086,-20641,-24334,-9828,6187,-23697),(280690,-30973,345,6263,12772,-38708,-23441,-14661,-9110,10692,13080,2834,8017,-7618,-5315,-3617),(291786,-32471,3395,5524,11964,-46644,-35581,-5547,-6530,10651,7272,-6194,16146,-2724,3191,4110),(263372,69779,8088,-26598,2552,-68406,-41601,1035,-22340,26423,-13963,14632,15588,-1813,-13939,-11868),(287536,-39043,-5308,10140,16379,-49009,-36987,-7954,-12075,16760,5980,-481,18783,148,-2853,2551),(291480,-39075,4110,6508,18038,-44824,-35765,-6204,-11397,11604,2636,-3210,13760,-212,1085,2332),(230759,-89863,-31554,35950,13284,-6547,-9001,11547,4930,5312,6215,-14609,3629,3279,2356,-6809),(291784,-42768,-1024,9570,19460,-43834,-33587,-8186,-12646,12821,4265,-1139,11335,-2055,-3220,-2158),(288903,-26613,-11381,5808,1421,-24756,-5776,-55629,-17211,24801,22582,36249,41501,9273,-19479,16296),(274485,-19209,-2363,3430,8804,-54436,-37994,-11056,-10936,20724,16464,1950,24739,7224,1281,8765),(222391,64518,-154902,37841,-26190,26823,-3123,-649,11992,-14394,-7319,-12479,-11563,-5018,938,-8888),(203601,85081,-144982,28034,-30830,24647,-452,-6440,12571,-15994,3894,-12425,-6213,-7693,-1203,-1065),(213239,114685,-140522,16459,-47099,34720,13306,-32802,14782,-20106,12828,-466,9220,-605,-4021,12319),(163322,110155,-94145,1548,-20096,-2360,-11870,-1856,-783,-799,-16987,7683,-11033,-9238,-13749,-15065),(218498,93806,-163701,31151,-40755,45470,14232,-28021,17614,-22308,10582,-1395,-132,-1672,-2646,9484),(216946,102433,-150913,24064,-42183,36915,12191,-30961,15666,-21656,15557,-1747,4289,-2886,-2860,13909),(159198,1743,-123025,44716,-19562,35144,8278,7728,19272,-10098,-245,-16798,-6822,-2370,3006,-63),(208440,71712,-118452,22154,-26971,4238,-10968,-15130,2391,-9705,9274,-14951,5001,679,1383,4458),(215276,97710,-135995,17968,-44886,63142,39362,-59206,14291,-19865,20131,28772,-3516,-4844,-16593,13587),(221217,83690,-144337,27595,-36441,22802,1777,-27147,10533,-13711,9151,-6773,6954,1148,524,9090),(325097,16968,-16193,-3112,-4904,20542,4515,25574,11770,-16943,-25152,-12600,-23068,269,6208,-14910),(268303,7500,38509,-20736,-4629,12465,14358,-4557,6818,-10594,-2474,2169,-10750,-2839,2650,1125),(275520,38185,32237,-26609,-20799,43022,41024,-21039,16779,-36507,14213,-9122,-23791,-11915,12247,4254),(265914,124449,33855,-54140,-27382,-11182,12505,-24711,-7301,7323,-2241,26120,8039,5667,-16793,1680),(251869,30333,34599,-24850,-12041,13576,16398,-104,12943,-18109,9301,-9232,-15380,-7727,8668,1689),(251869,30333,34599,-24850,-12041,13576,16398,-104,12943,-18109,9301,-9232,-15380,-7727,8668,1689),(325989,-57911,-30082,21851,-6573,45563,24684,29129,23692,-6355,-28650,-2923,-327,10845,3034,5258),(280155,37672,52645,-35777,-19963,12117,14858,1461,14287,-8099,5226,-9650,5493,7484,14025,19528),(276828,10302,52179,-29632,-15267,39793,47098,-52080,-5453,-9639,10309,31347,9921,12898,-8657,13019),(260791,23896,44968,-26734,-4326,-1042,-2253,18580,9705,-16199,-12736,-21284,-12144,747,16458,-1234),(214135,-62139,-11501,19982,16803,-22738,-8962,6822,-13691,18468,-3655,14301,673,-2218,-15760,-23495),(270812,-37830,143,8886,13546,-43327,-30336,11202,-19837,16938,188,-2322,2937,-4406,-9326,-13584),(276217,-38499,11308,4297,9673,-47861,-28956,7183,-16177,22889,3332,1799,16414,-3452,-11546,-1344),(165659,47466,32763,-27428,-205,-51973,-27846,10064,-16421,19924,-2475,3944,5265,5,-2100,-12757),(266082,-33761,7985,4878,12729,-40541,-32175,13648,-15489,12581,3172,-10668,-80,-4188,-1920,-11375),(254210,-52366,-5196,14975,16730,-35175,-21368,6553,-19136,18164,-2859,6504,-258,-4661,-16105,-19144),(127837,-75797,-36620,34532,11309,7025,3782,5062,-991,4040,901,3606,-3261,-3286,-12483,-11031),(269700,-38604,16353,3102,13444,-44926,-28783,13963,-15341,14326,4675,-9796,4366,-6409,-5387,-8712),(265314,-31109,-356,5227,500,-47960,-25272,-7863,-16641,38652,15327,16852,37194,7952,-17538,15990),(259177,-38887,7442,6560,13703,-41392,-25285,12124,-16911,16715,-2052,-1886,706,-7522,-10000,-14983),(292046,-37559,-37454,20933,6676,-24300,-19387,14671,-4530,21394,-12696,6528,14417,6219,-9207,-12707),(262416,-21513,-16840,9952,1230,-39882,-28923,11256,-1204,22369,9708,-1883,17931,4512,655,7452),(291716,-10524,-39086,14943,-2942,-39053,-31447,391,-1483,15553,14920,-2889,22086,3795,3014,9920),(236642,85409,9038,-31280,-11220,-46438,-28472,20020,-7497,22409,-16732,3234,8422,4653,-210,-6498),(281347,-1069,-33074,10696,-3661,-34522,-32389,13232,1448,7134,12909,-16582,10628,2655,12556,8260),(281347,-1069,-33074,10696,-3661,-34522,-32389,13232,1448,7134,12909,-16582,10628,2655,12556,8260),(189039,-80821,-57864,42872,3670,30878,13788,18040,14252,-3406,-6474,-5807,-8234,182,-931,-2524),(272788,-19914,-30842,15029,4305,-43367,-36867,6333,-6505,17848,12827,-4836,15175,2829,3966,5220),(269795,-4935,-31350,10512,-6561,-33171,-25098,-9191,-1046,13667,28663,-2289,19582,5844,1457,15022),(282694,12486,-26722,2258,-18913,-28289,-16401,-9019,1665,18900,30703,4828,35736,10245,4604,28754),(246490,-40028,-10131,12617,7452,7212,3458,3102,-3972,-3399,-6239,3192,-11652,-2662,-1479,-13537),(317755,-47367,47566,-9880,8103,33620,29091,-79,-3068,-16491,-18458,16332,-16874,-6220,1560,-6989),(334261,-19166,42226,-13663,3296,21948,9363,30359,9341,-33161,-23471,-22231,-30456,-12213,23132,-11694),(184795,72766,29784,-34131,-6333,-32692,-19590,21383,-5303,9230,-13409,-2954,-7180,-160,7454,-13493),(344569,-16602,38324,-15646,-5530,30066,19239,-309,721,-18642,-10178,5070,-6995,-5528,12142,9244),(341190,-16990,21464,-5872,6021,26322,6947,32040,9512,-37394,-19978,-28718,-42999,-19283,24077,-17899),(214015,-99966,-59776,48281,2794,66941,34769,20390,21975,-22393,-15374,-9495,-20217,-3444,4211,-865),(326484,-13597,30179,-9535,9071,10824,-3469,38722,7343,-29076,-15711,-33385,-44010,-16713,26856,-20484),(329638,-36502,29642,-6490,4213,30935,21006,-14340,-11146,-19253,-8497,19030,-10050,-5155,7699,543),(314798,2635,25747,-13539,-6756,7062,943,32153,11655,-17744,-5965,-19463,-17387,-5770,22588,876));
			w_2D := ((44,28,17,9,7,7,10,14,16,18,20,20,21,22,23,24,25,27,28,28,26,23,20,17,14,10,7,7,9,12,21,33,39,22,10,7,6,10,15,18,21,24,26,29,30,31,32,33,34,35,34,35,32,28,24,20,17,13,8,6,7,10,16,28,32,17,8,5,8,13,18,21,23,27,32,35,36,37,37,38,38,38,38,38,36,31,26,23,20,15,11,6,5,8,14,25,28,12,5,6,10,16,21,23,25,29,33,36,39,40,40,40,40,40,39,39,36,32,28,25,22,18,13,7,5,6,12,22,26,8,5,6,12,18,22,25,27,30,34,38,41,42,42,41,41,41,40,39,36,33,29,26,23,19,14,8,4,4,10,19,23,6,4,6,13,19,23,27,29,33,36,41,43,43,43,43,43,42,42,41,38,33,29,27,24,21,15,9,4,4,9,17,20,6,4,6,14,20,24,28,31,35,40,44,46,45,45,44,45,44,44,43,39,35,30,27,24,21,17,10,5,3,8,17,19,5,4,7,16,22,25,28,31,35,39,42,44,45,46,46,46,45,42,40,36,32,29,26,24,22,19,12,6,3,7,15,18,5,4,8,19,24,25,22,22,23,26,30,33,38,41,43,41,37,32,26,23,20,18,18,20,21,21,15,8,4,8,16,18,6,4,10,21,24,19,16,16,13,13,16,20,25,31,35,33,27,19,14,13,13,14,14,14,17,19,17,11,5,8,14,19,6,5,12,23,21,17,17,19,17,14,13,13,17,25,31,28,20,15,13,14,17,18,18,17,17,19,19,13,6,8,14,22,8,7,15,22,22,20,19,18,19,16,14,14,16,24,34,31,20,14,14,15,16,18,16,17,19,21,21,16,8,9,15,26,11,8,17,25,25,22,16,15,11,8,12,13,15,24,40,41,24,14,13,13,9,10,13,15,20,23,23,19,10,10,17,31,16,10,20,29,28,22,17,19,15,13,18,16,21,26,43,45,27,21,17,18,15,17,19,19,22,25,26,22,14,13,20,36,22,15,23,31,31,28,25,22,22,21,21,24,28,30,44,47,29,27,24,20,21,22,23,26,28,29,29,24,17,15,22,40,24,18,24,33,33,34,33,31,29,28,30,35,31,33,45,49,32,28,33,32,30,32,34,34,34,32,29,26,18,17,25,44,26,21,24,33,35,37,39,40,40,39,41,37,30,34,46,51,35,29,32,38,39,39,40,40,37,33,30,27,20,20,29,49,32,25,25,33,35,38,42,44,42,44,42,33,30,36,47,51,37,29,28,37,41,41,41,39,35,31,29,26,21,23,32,53,39,28,26,31,33,36,39,42,42,42,38,30,33,36,45,48,35,30,27,31,37,39,38,35,32,29,29,27,24,29,35,57,43,33,28,30,31,33,36,39,40,38,34,30,32,30,35,36,29,27,27,26,31,35,34,32,30,28,26,26,27,31,38,58,48,36,30,29,30,31,33,35,37,35,31,27,19,18,23,24,20,18,22,26,27,30,30,29,27,25,25,25,28,35,43,60,54,42,35,29,29,29,29,32,32,31,30,26,19,14,16,16,15,14,22,27,27,26,26,26,25,24,25,28,31,40,49,62,60,50,40,30,27,27,27,29,29,29,28,26,22,21,18,17,18,19,22,24,26,25,24,24,23,23,25,31,39,48,53,64,63,56,46,33,27,26,26,26,26,25,24,23,21,22,22,22,21,21,20,20,20,22,23,24,23,22,26,34,44,51,57,64,63,60,53,40,27,25,25,26,24,21,18,16,17,17,18,20,17,16,15,15,16,19,23,24,22,23,29,40,49,55,58,65,63,62,58,46,30,25,25,25,23,19,15,15,14,16,18,17,17,15,14,14,16,18,22,24,22,23,32,43,52,57,60,65,64,63,59,51,33,26,25,24,23,19,19,19,17,19,21,20,20,18,17,19,19,19,21,22,21,26,37,47,55,59,61,66,65,64,61,55,38,27,25,23,22,21,22,22,20,18,17,16,17,18,19,21,21,20,20,20,22,29,41,51,59,61,61,66,65,65,64,58,44,29,24,22,21,22,23,23,22,21,20,20,21,21,22,22,21,20,20,19,22,31,43,51,59,61,61,68,67,65,64,59,48,35,23,21,20,22,24,25,25,26,28,28,28,28,26,24,22,20,19,18,22,32,43,54,58,59,60,68,67,66,65,58,47,37,26,20,19,20,23,25,26,28,29,28,28,27,25,23,21,18,16,18,22,31,39,51,55,57,60,67,67,66,63,54,43,37,25,19,18,18,19,22,24,25,24,24,22,22,21,19,18,16,15,17,22,29,36,45,54,57,59),(31,41,46,34,25,15,17,26,34,32,30,29,27,26,23,18,12,4,-2,-6,-9,-9,-9,-6,-1,0,10,11,11,12,2,-27,35,50,33,26,13,12,23,32,32,32,28,25,22,18,13,8,0,-6,-11,-16,-19,-19,-17,-14,-8,-3,0,5,10,9,3,-18,46,49,29,14,8,18,28,30,32,30,26,24,16,11,3,-2,-8,-14,-17,-22,-26,-26,-23,-20,-15,-9,-5,0,5,8,0,-19,46,36,16,11,8,21,27,28,29,28,27,19,12,4,-3,-10,-15,-17,-18,-23,-26,-27,-26,-25,-22,-15,-10,-4,0,2,-3,-19,47,27,15,8,11,22,27,27,28,28,22,15,7,-2,-11,-14,-17,-18,-19,-25,-27,-28,-28,-29,-27,-21,-15,-8,-2,0,-3,-17,38,17,12,9,13,22,26,25,25,23,16,11,2,-10,-16,-17,-19,-20,-22,-27,-29,-30,-30,-30,-29,-26,-20,-11,-4,-1,-3,-13,25,15,11,9,13,19,22,22,20,17,12,6,-3,-14,-19,-22,-22,-22,-25,-30,-33,-32,-31,-31,-30,-27,-23,-14,-9,-2,-3,-19,18,13,10,8,11,18,21,17,16,15,11,4,-7,-13,-17,-19,-20,-20,-22,-27,-29,-30,-29,-27,-27,-28,-26,-19,-13,-5,-7,-23,14,12,9,6,8,20,26,27,27,28,24,13,7,0,-4,-4,-11,-11,-12,-13,-12,-8,-5,-5,-13,-20,-24,-23,-15,-6,-10,-27,8,11,8,3,8,23,37,31,26,20,12,10,16,18,18,15,4,0,-2,2,10,9,6,0,-2,-6,-18,-22,-18,-7,-10,-27,14,11,7,0,11,28,34,31,14,13,10,12,20,26,34,34,13,-1,-2,3,8,5,0,-5,-7,-9,-12,-17,-16,-7,-14,-31,11,11,1,2,19,32,32,23,14,0,-8,1,10,25,43,47,24,-5,-9,-1,0,-3,-13,-13,-14,-15,-17,-14,-15,-10,-23,-37,14,8,2,0,23,36,34,24,20,8,0,9,10,20,40,41,18,-9,-11,-1,7,14,-3,-4,-5,-13,-15,-15,-14,-12,-25,-43,17,8,2,2,27,42,35,30,27,19,12,9,17,20,37,35,9,-6,-6,1,7,18,6,-1,0,-7,-12,-16,-11,-18,-29,-49,17,14,1,6,34,42,41,39,37,35,34,30,30,36,39,29,3,-9,-2,6,8,12,12,9,0,-3,-9,-18,-17,-23,-38,-55,22,17,3,6,36,43,43,44,50,53,45,41,41,36,39,28,0,-10,-6,-2,12,17,17,14,8,1,-9,-15,-19,-24,-43,-65,20,18,12,7,35,42,44,45,45,46,44,45,37,42,38,28,-2,-11,-11,-9,0,7,12,8,1,-7,-14,-18,-24,-30,-47,-77,16,14,11,7,36,40,41,41,43,46,44,44,42,38,36,27,-3,-17,-14,-12,-7,-1,2,1,-6,-13,-19,-23,-27,-35,-54,-81,10,13,6,9,35,40,41,41,46,47,47,44,41,32,25,19,-10,-23,-15,-19,-10,0,0,-2,-8,-16,-22,-26,-29,-45,-71,-79,4,14,10,13,32,42,42,41,44,48,47,43,31,19,9,4,-15,-30,-23,-19,-10,-6,0,-4,-12,-20,-24,-24,-31,-50,-72,-86,2,12,12,16,29,41,42,42,44,44,40,37,30,19,17,12,-4,-18,-24,-9,-4,-2,0,-5,-14,-20,-22,-24,-34,-54,-79,-92,1,3,10,14,28,40,40,40,42,41,37,39,39,30,27,18,7,7,6,2,-4,0,-2,-7,-14,-19,-21,-27,-38,-62,-89,-94,-5,-6,6,15,26,38,41,41,43,42,38,36,35,36,33,21,16,17,12,5,-3,-4,0,-9,-15,-17,-21,-31,-51,-75,-90,-97,-9,-13,-3,17,24,35,41,41,42,39,35,36,38,36,34,29,24,16,11,5,-1,-2,0,-6,-14,-16,-20,-37,-56,-86,-94,-94,-9,-12,-9,0,20,34,41,42,42,35,30,32,30,27,24,18,13,6,1,-1,-3,-3,-2,-4,-9,-16,-22,-46,-76,-94,-95,-92,-5,-12,-8,-2,12,34,43,46,46,35,28,22,20,15,10,3,2,0,-4,-9,-8,-4,-2,-2,-8,-15,-25,-54,-87,-97,-94,-88,-4,-11,-12,-7,9,32,41,48,50,42,33,32,32,27,24,16,11,6,2,-1,-2,0,3,-1,-8,-13,-35,-66,-94,-95,-85,-80,-3,-8,-11,-8,3,25,39,45,49,48,41,42,42,36,26,21,17,13,8,2,2,3,3,-1,-8,-17,-46,-81,-96,-90,-78,-78,6,1,-1,-3,3,16,39,45,49,45,42,43,42,35,28,27,25,24,20,10,5,3,2,-1,-7,-25,-56,-84,-91,-79,-71,-67,15,8,11,5,18,26,33,50,47,46,44,43,42,39,38,34,29,26,20,13,8,3,1,-1,-8,-31,-62,-81,-88,-82,-76,-76,23,23,22,21,27,34,36,43,48,46,46,44,46,47,46,39,36,30,21,13,7,3,0,-2,-15,-35,-60,-75,-77,-88,-82,-74,26,35,33,32,34,44,41,40,43,42,43,45,45,45,43,36,35,31,22,13,5,1,0,-6,-22,-40,-51,-62,-67,-84,-88,-82),(7,18,26,6,3,-2,8,20,25,32,38,40,40,43,46,48,47,48,46,42,32,21,13,10,4,1,6,10,18,29,40,34,15,21,9,6,0,9,25,31,37,43,46,49,50,51,50,52,51,48,47,45,37,26,16,10,6,2,3,7,11,22,29,39,26,24,4,2,5,23,34,38,42,45,51,51,50,51,50,50,48,45,46,43,35,25,19,14,8,3,2,4,6,16,32,33,27,21,7,3,11,30,38,40,42,44,48,47,44,47,48,47,45,43,42,37,31,23,19,16,12,7,3,3,4,9,30,31,38,10,5,7,16,32,38,41,41,42,45,45,41,46,48,48,47,45,42,37,32,24,20,16,13,7,5,2,0,5,22,35,39,9,5,8,20,33,38,41,42,42,42,39,39,49,52,50,49,48,46,42,34,24,21,17,14,8,5,2,-1,2,17,35,37,10,5,9,21,35,39,40,41,37,35,35,44,49,50,49,49,45,44,37,29,23,21,17,14,8,6,3,-1,0,14,30,37,11,6,10,23,35,36,36,31,26,27,32,40,41,42,45,43,39,33,27,21,19,17,16,12,5,5,5,-2,0,9,22,44,10,7,12,27,33,26,17,10,7,12,19,21,22,23,22,18,17,10,4,0,-4,-5,-6,0,-1,3,6,-2,-2,8,18,47,13,8,13,25,22,0,-24,-23,-23,-16,-14,-15,-10,-8,-8,-15,-17,-24,-24,-30,-31,-31,-32,-30,-21,-6,4,-1,-3,7,12,50,16,8,13,21,7,-27,-32,-26,-30,-32,-27,-24,-22,-23,-26,-38,-39,-35,-28,-24,-26,-23,-26,-35,-37,-22,-8,-9,-8,3,13,56,24,11,9,15,-4,-17,-9,-3,-5,-11,-21,-21,-19,-25,-35,-50,-42,-26,-17,-18,-16,-10,-17,-19,-27,-26,-18,-12,-11,0,16,57,28,11,8,10,-5,-1,-5,-9,2,-10,-19,-18,-19,-28,-38,-48,-38,-29,-23,-22,-20,-17,-27,-27,-32,-34,-29,-18,-14,0,16,59,40,17,11,7,-9,-12,-19,-19,-21,-27,-22,-30,-25,-24,-29,-38,-41,-40,-34,-33,-39,-40,-45,-45,-41,-40,-32,-22,-17,2,15,61,43,24,14,3,-15,-22,-24,-30,-28,-32,-35,-37,-33,-23,-28,-37,-38,-46,-53,-49,-47,-53,-58,-50,-45,-41,-34,-27,-18,0,9,57,32,27,11,-2,-17,-26,-34,-39,-42,-39,-41,-27,-28,-21,-28,-32,-40,-47,-42,-52,-53,-49,-48,-51,-50,-42,-35,-28,-17,1,1,54,35,27,9,-8,-15,-27,-32,-30,-30,-28,-26,-19,-25,-19,-24,-26,-36,-42,-44,-44,-48,-47,-44,-48,-43,-40,-33,-27,-13,0,-2,56,39,27,9,-2,-9,-18,-26,-26,-27,-24,-22,-18,-19,-18,-22,-26,-31,-39,-38,-42,-44,-43,-41,-42,-40,-37,-32,-24,-10,-6,2,57,50,30,17,4,-9,-12,-17,-26,-26,-23,-21,-16,-19,-15,-11,-21,-30,-40,-30,-41,-47,-43,-41,-41,-39,-35,-30,-22,-6,-4,1,55,48,45,28,10,-4,-11,-16,-22,-25,-21,-22,-15,-10,-7,-9,-14,-21,-28,-30,-34,-37,-42,-43,-40,-34,-31,-28,-23,-5,-5,-2,53,48,44,33,14,0,-8,-12,-16,-22,-27,-23,-15,-4,-2,-7,-13,-15,-20,-37,-48,-35,-36,-39,-37,-33,-30,-27,-20,-7,-5,4,52,49,46,41,20,3,-6,-12,-17,-22,-29,-28,-20,-12,-20,-19,-23,-31,-39,-42,-45,-48,-36,-32,-34,-32,-28,-24,-19,-14,-2,2,52,51,46,46,27,6,-5,-11,-18,-26,-30,-28,-30,-38,-40,-39,-38,-49,-52,-50,-48,-47,-44,-35,-32,-31,-27,-21,-18,-7,7,9,53,53,53,52,35,9,-2,-9,-14,-22,-29,-32,-36,-40,-43,-46,-44,-46,-48,-49,-47,-45,-43,-40,-35,-31,-28,-23,-9,-1,8,10,47,52,54,58,46,13,-1,-7,-12,-23,-27,-25,-23,-25,-28,-28,-30,-25,-30,-32,-31,-30,-35,-41,-40,-33,-29,-22,-7,3,10,12,37,50,56,63,54,26,0,-9,-17,-25,-22,-15,-10,-6,-5,-8,-11,-14,-15,-19,-23,-24,-30,-42,-43,-34,-29,-17,-2,3,11,12,36,51,57,60,59,36,2,-12,-21,-27,-20,-9,-5,-10,-12,-15,-18,-20,-27,-34,-36,-37,-34,-40,-41,-36,-29,-16,4,5,-4,-12,33,44,48,55,62,49,12,-11,-18,-24,-27,-21,-18,-17,-20,-21,-23,-29,-35,-40,-42,-41,-41,-38,-37,-35,-29,-8,-1,-8,-15,-17,17,28,35,41,56,48,20,-5,-16,-20,-26,-23,-20,-21,-29,-40,-49,-52,-51,-46,-42,-42,-42,-40,-38,-38,-31,-15,-13,-28,-27,-34,1,12,23,36,36,24,16,-9,-16,-19,-23,-24,-25,-30,-35,-41,-44,-48,-48,-46,-46,-43,-42,-42,-40,-43,-35,-26,-15,-21,-19,-19,-9,4,11,18,12,0,6,-3,-15,-21,-25,-28,-31,-39,-40,-40,-43,-45,-51,-53,-50,-45,-42,-38,-37,-42,-41,-34,-23,-17,-19,-20,-6,2,4,9,-6,-12,-3,0,-8,-17,-26,-29,-30,-34,-34,-36,-43,-48,-50,-50,-46,-41,-37,-31,-31,-39,-40,-44,-30,-14,-14,-6),(-17,-24,-29,-12,-10,-5,-8,-13,-20,-21,-23,-23,-22,-26,-26,-25,-24,-20,-17,-12,-10,-3,-2,-2,1,0,-6,-7,-12,-16,-19,-11,-24,-30,-16,-10,-2,-7,-17,-20,-24,-25,-27,-26,-23,-24,-24,-23,-18,-16,-16,-13,-8,-6,0,3,2,2,0,-2,-8,-12,-17,-17,-29,-31,-13,-6,-3,-12,-21,-22,-25,-27,-26,-24,-24,-21,-21,-19,-17,-14,-12,-9,-4,-3,-2,0,0,2,1,-3,-5,-9,-14,-12,-31,-22,-7,-3,-6,-17,-23,-23,-23,-24,-27,-21,-18,-18,-17,-16,-12,-10,-9,-8,-4,0,0,0,2,2,4,0,-2,-6,-14,-9,-34,-12,-7,-4,-9,-18,-23,-22,-23,-25,-23,-19,-18,-14,-11,-13,-14,-12,-10,-7,-4,-1,0,0,1,3,5,3,0,0,-7,-11,-33,-10,-5,-5,-9,-17,-21,-21,-20,-22,-18,-18,-15,-12,-14,-12,-12,-12,-9,-5,-5,1,0,2,2,4,5,3,2,-1,-7,-13,-26,-9,-5,-6,-11,-18,-21,-20,-19,-17,-15,-12,-12,-11,-13,-12,-12,-9,-8,-4,-1,3,2,1,1,3,4,4,3,0,-6,-6,-21,-7,-6,-7,-13,-19,-19,-17,-15,-13,-12,-12,-12,-10,-9,-9,-10,-6,-5,0,0,0,3,1,1,8,6,4,5,2,-1,-3,-25,-5,-6,-4,-12,-16,-17,-13,-10,-9,-11,-12,-8,-7,-7,-4,-4,-2,4,3,8,7,4,4,2,7,5,2,5,1,1,0,-21,-10,-8,-3,-10,-15,-10,0,2,1,2,2,0,0,0,0,5,6,9,8,9,10,10,10,9,7,6,6,8,6,1,2,-26,-10,-3,-6,-8,-11,2,1,2,7,6,8,2,1,-1,-1,12,18,16,9,8,7,11,9,17,16,11,10,10,4,4,1,-27,-13,-5,-4,-8,-5,-2,-1,-3,1,7,7,4,0,-5,1,13,17,13,6,5,5,7,10,13,15,15,12,8,9,6,0,-32,-15,-5,-3,-9,-8,-10,-6,-3,-3,5,5,4,1,-3,1,15,20,11,8,4,5,7,9,12,17,16,17,13,8,5,2,-30,-19,-8,-5,-11,-8,-4,-2,-1,3,5,5,3,3,0,-1,12,18,17,12,11,12,14,18,16,16,16,17,14,12,6,5,-31,-24,-11,-4,-12,-8,-2,-1,0,1,1,3,5,2,-2,3,15,16,18,19,14,14,14,17,15,18,18,19,15,14,7,7,-32,-18,-12,-5,-8,-6,-1,1,0,1,0,2,-1,1,-5,0,13,21,17,17,16,15,12,11,17,20,18,16,17,12,10,13,-32,-24,-15,-4,-9,-8,-4,0,-2,0,-2,-2,-3,-1,-4,0,11,17,20,19,17,18,15,15,17,19,21,19,16,12,11,15,-32,-23,-15,-5,-10,-7,-6,-3,-1,-2,-2,-3,-6,-2,-4,0,12,16,20,16,18,17,16,14,18,21,18,20,17,13,14,14,-27,-28,-15,-11,-10,-8,-8,-7,-2,-4,-4,-4,-5,-4,0,-1,12,19,20,16,16,17,16,15,21,19,19,20,16,12,14,18,-25,-27,-22,-14,-12,-10,-6,-6,-3,-3,-6,-3,-1,-1,-1,2,11,17,18,15,13,13,15,17,19,19,17,16,15,12,15,19,-24,-27,-22,-18,-14,-12,-9,-6,-5,-6,-2,-3,-1,-3,-4,-2,8,11,14,16,19,14,12,15,16,16,18,17,16,15,20,21,-22,-23,-25,-22,-17,-14,-12,-9,-6,-6,-1,-1,-6,-6,0,2,4,8,9,12,16,16,12,13,16,16,17,14,14,18,24,24,-19,-19,-20,-23,-20,-16,-11,-10,-6,-2,0,-2,1,1,4,8,8,10,14,14,18,18,15,15,17,17,17,14,16,19,19,22,-18,-17,-21,-26,-23,-17,-13,-10,-8,-4,-1,0,1,2,7,8,8,11,14,13,17,17,16,14,16,16,15,15,15,21,20,24,-15,-15,-20,-26,-27,-17,-11,-10,-8,-4,1,-1,0,1,1,5,8,5,10,11,12,10,12,15,18,17,16,19,20,22,22,22,-9,-15,-17,-27,-28,-24,-13,-12,-10,-3,-1,-2,-2,-2,0,4,4,6,7,10,10,12,9,15,19,17,14,17,21,25,21,21,-11,-16,-17,-22,-28,-29,-16,-9,-9,-3,-1,-5,-7,-3,-2,3,4,7,10,13,15,10,11,16,17,15,18,18,23,24,27,29,-10,-13,-13,-18,-26,-30,-22,-11,-7,-6,-2,-5,-5,-3,1,2,3,5,9,14,12,12,16,14,16,16,18,22,25,28,30,29,-6,-9,-9,-13,-22,-24,-24,-13,-9,-7,-4,-2,-4,-5,0,5,8,11,12,11,12,15,13,16,17,19,24,30,34,36,32,33,-3,-6,-9,-13,-18,-19,-18,-15,-9,-7,-6,-4,-4,-1,0,5,8,10,12,13,16,15,16,13,15,21,30,36,32,32,31,31,-3,-5,-10,-10,-7,-6,-16,-14,-8,-7,-4,-4,-1,3,3,5,7,9,15,15,16,14,16,13,15,22,32,35,32,34,33,29,-3,-10,-7,-7,-3,-5,-8,-11,-9,-5,-2,-2,-1,0,2,2,6,9,11,13,13,15,13,12,16,22,26,36,34,34,33,29),(-39,-49,-45,-27,-15,0,-5,-2,1,-11,-1,4,-7,0,-2,-4,-3,-13,-12,-1,-1,-8,-9,-10,-12,-8,-6,-8,-7,-22,-28,-24,-50,-61,-28,-16,-8,6,-4,-2,-10,-10,-2,8,-7,-11,3,2,-4,2,0,0,0,1,-14,-8,-16,-14,-8,-16,-13,-11,-8,-16,-66,-43,-13,-1,-9,-13,-3,-8,-1,7,0,4,2,-4,2,3,12,10,11,12,0,3,0,-6,4,-11,-11,-4,0,-14,-12,-24,-59,-43,-20,-2,-2,2,-10,-2,2,-7,2,3,-3,4,18,12,16,3,4,5,-5,-6,1,-2,-7,-10,-2,-6,2,-5,0,-8,-64,-29,1,-5,8,-1,0,-2,-1,5,5,1,6,3,7,7,14,11,9,-1,-2,5,5,-3,0,0,-12,-4,0,-2,-6,0,-54,-17,-3,3,-2,-8,8,1,-1,6,8,17,9,0,12,10,17,15,11,7,13,-1,9,5,-3,-6,-12,-4,-2,-4,-2,-5,-45,-5,-8,1,-5,0,13,9,10,11,8,3,6,6,16,24,9,16,7,13,8,-1,-2,-3,-2,-2,-3,-10,-1,-7,5,1,-39,-21,-7,-9,3,6,-4,6,5,15,17,15,20,22,19,12,11,16,24,10,17,9,-6,-1,0,-1,-7,1,3,-6,-3,-6,-22,-16,3,-11,12,7,0,7,5,5,14,20,10,7,8,4,23,4,2,19,0,-3,-2,2,1,-12,-3,0,3,-1,-3,5,-34,0,0,-4,6,9,0,-2,0,5,0,3,6,8,-3,-12,0,2,4,11,0,-5,0,1,3,0,-12,0,-4,-11,-9,13,-39,-11,-8,12,7,7,3,-1,10,-11,-5,-11,0,-3,-17,-10,-8,-6,-7,-9,-6,6,-6,-7,-14,-14,-14,-4,-5,0,-8,11,-31,-9,-1,12,15,-13,-9,-10,5,6,2,-9,0,2,-5,-12,-3,6,2,6,-3,2,12,-7,-4,-5,5,-10,-2,-10,3,9,-37,-14,-2,14,16,-3,0,-4,6,-10,-12,10,-10,-1,3,2,4,-9,-6,1,2,2,-3,-5,-11,-18,-4,-5,-13,-1,-3,13,-38,-9,8,13,12,3,-1,-1,14,1,13,9,-1,8,-14,-1,5,-12,-9,-8,0,-11,-5,-10,2,-3,-8,-12,-3,-3,4,1,-26,-7,-4,6,14,-12,-14,-12,-10,-4,-3,0,-5,-1,0,12,-2,2,-17,-13,-1,-12,3,-5,-15,-6,-7,-4,-11,-8,7,15,-25,-16,-7,0,-1,3,-8,-9,-10,-4,-8,0,-4,-3,9,-3,7,-5,-6,-9,-15,-10,-11,-21,-21,-14,-1,0,-12,-2,11,17,-7,-11,-9,11,-2,-3,-7,-3,0,-6,2,0,2,-1,-7,0,6,0,-4,-11,-19,-12,-18,-18,-8,-9,-6,-7,-8,0,23,26,-1,-15,-10,2,5,-3,-4,-1,-4,3,-9,-6,0,-15,-8,-4,-4,8,-1,-5,-16,-12,-6,1,-6,-8,-5,-4,-3,-4,19,29,1,-14,-10,3,-6,-2,-6,3,-1,-9,-10,3,-12,5,-2,4,13,-5,-8,4,-8,-12,-8,2,-12,-4,0,-5,-11,6,20,25,10,0,-12,-3,-6,-7,-4,-3,4,2,-5,-2,1,3,4,4,11,-6,-2,0,5,-1,-5,-5,-2,-5,-1,-5,2,5,25,22,8,3,-7,-16,-7,8,-5,-3,0,1,0,-6,0,5,-3,5,4,8,-2,0,-1,-3,0,-3,-2,-7,-3,-4,-8,2,27,29,3,3,7,-8,-18,6,3,-1,-4,6,-1,-3,0,-6,-6,6,5,2,-1,-11,-8,0,-4,-4,-9,-5,-7,-10,6,8,28,32,12,3,0,5,-20,3,2,6,-7,0,-5,-2,-4,0,-12,4,1,1,-9,-2,-6,-7,-9,-4,-5,-12,-6,3,0,20,33,35,17,17,10,-5,-17,-14,-10,10,1,2,2,9,0,2,-4,-12,-13,-5,-18,-1,-1,-4,-9,-18,-5,-14,0,-2,9,22,36,25,22,16,18,-4,-17,-4,-2,4,-9,-4,-3,-2,0,-7,5,-11,-9,-2,9,-6,1,-4,-6,-1,-6,-11,-7,-1,15,31,21,13,2,9,4,7,-16,-19,-14,3,-6,-3,0,-2,8,7,-2,-5,12,9,-9,-10,-10,-9,0,-3,-16,-3,-14,1,28,34,15,18,10,13,13,6,-1,-19,-5,-13,-2,-1,-9,-6,-12,-3,4,0,-1,-1,2,-5,-14,-6,-5,-16,-3,-2,-15,19,23,25,17,18,14,14,8,13,-11,-18,-6,-2,-14,-3,5,-3,-2,-8,-3,-10,-4,0,-6,-11,-3,-14,-11,-17,-6,-10,0,24,28,16,12,11,4,13,3,10,-6,-14,-28,-19,-13,-10,-13,-11,-6,-5,-11,-15,0,-19,-17,-15,-17,-9,-12,-20,-18,-6,7,25,13,10,9,3,-4,-3,-4,-3,-14,-5,-22,-13,-16,-15,-14,-10,-12,-18,-6,-16,-9,-21,-11,-12,-21,-22,-16,-4,-21,-13,10,22,12,23,19,11,-5,2,3,-2,-15,-14,-14,-9,-22,-21,-4,-1,-19,-19,-26,-24,-25,-19,-18,-12,-12,-23,-13,-2,-1,-1,7,18,13,14,14,10,-7,6,-8,-5,7,-13,-15,-12,-19,-19,-13,1,1,-6,-14,-8,-14,-28,-16,-14,-6,-11,-7,-12,0,4,8,5,15,11,19,12),(9,39,58,31,35,24,33,31,52,51,43,34,47,57,54,54,64,48,64,37,46,38,40,46,39,38,45,52,61,84,88,91,38,53,37,24,6,32,40,44,52,49,53,40,46,52,35,42,36,37,45,42,33,40,40,35,45,40,41,44,53,67,93,104,49,45,34,25,17,28,41,38,40,44,42,24,37,30,36,26,23,28,21,20,24,30,44,48,46,36,26,38,44,60,72,112,50,44,20,10,25,35,53,42,29,34,31,15,15,24,-1,16,1,14,15,15,25,28,31,49,37,46,27,25,28,45,81,96,43,21,8,12,23,32,27,15,32,15,18,16,8,7,-4,0,1,2,17,15,26,16,35,47,35,32,26,17,19,27,61,85,52,28,20,16,23,26,12,9,8,12,-7,-5,-3,-11,-12,-8,-11,-3,-6,6,24,10,18,27,36,35,26,15,11,24,56,86,53,24,7,12,21,12,1,1,0,0,-6,-2,-22,-14,-10,-19,-3,-18,-7,5,6,2,19,28,39,35,27,25,13,20,47,78,35,15,15,17,10,3,-3,3,5,-3,-12,-7,-9,-17,-15,-18,-14,-34,-20,-9,-12,4,-2,18,31,23,29,23,11,5,29,76,41,11,16,0,-5,-14,5,5,14,8,1,-1,1,3,-8,-21,-15,-19,-19,-14,-14,-3,-5,2,13,22,35,33,13,24,28,68,34,17,23,-15,-14,-7,4,-6,-12,3,-7,-6,-1,-7,-9,-3,-5,-9,7,-4,0,0,12,6,16,24,39,21,8,13,34,54,44,19,13,-13,-31,-22,-25,-11,-23,-34,-18,-25,-18,-10,-6,15,9,-5,1,-4,-17,-12,-19,4,19,23,37,20,5,18,32,58,19,13,4,-21,-31,-16,-13,-27,-24,-23,-26,-18,-15,-19,-8,0,14,0,-11,-24,-22,-22,-18,3,-4,23,33,31,26,16,39,56,31,24,1,-25,-28,-19,-13,-11,-19,4,7,-15,-17,-18,-3,-1,3,-1,0,-16,-9,-14,0,19,11,22,37,28,28,30,41,49,22,13,0,-23,-21,-15,-22,-21,-31,-37,-40,-24,-4,-26,-10,0,4,8,19,-1,-9,-11,11,13,21,31,40,25,22,19,46,48,5,8,8,-29,-9,0,-13,-10,-5,-11,-5,-10,-15,-20,-17,-22,-11,26,26,12,22,15,9,35,43,31,32,15,25,19,46,47,-4,-6,-2,-20,-16,0,-11,-22,-11,-17,-2,-16,-7,-12,-17,-9,-8,6,22,20,26,26,23,41,33,30,20,24,40,27,30,38,-21,-3,-8,-43,-10,6,0,-6,6,-1,-11,-10,-7,-12,-20,-22,-5,4,21,29,37,15,22,35,27,12,20,23,33,28,15,32,-32,-11,-17,-39,-20,-12,0,0,-7,-7,-3,-11,3,-7,-13,-16,-9,1,15,18,31,24,12,15,15,5,30,21,25,23,22,14,-48,-9,-16,-24,-16,-13,-9,-5,-19,0,-4,1,-5,-22,-27,-22,-15,9,19,9,33,27,16,17,4,20,13,13,25,23,12,-12,-58,-53,-14,-27,-30,-10,-19,-9,-19,-3,0,-4,-29,-27,-14,-32,-21,1,-6,12,30,19,22,11,11,13,25,30,13,6,6,2,-53,-58,-34,-17,-16,-13,-17,-17,-13,-1,-9,-1,-20,-20,-28,-26,-13,-3,1,16,15,16,20,10,18,29,18,23,9,-1,-2,-6,-54,-52,-41,-24,-16,-16,-10,-1,-10,-4,-17,0,10,10,-12,-19,1,19,29,33,20,12,16,21,23,18,18,29,22,6,-25,-14,-58,-58,-59,-26,-9,-4,-9,-6,-3,-16,-14,8,-12,2,7,1,-4,18,26,16,14,20,24,18,16,20,27,25,22,24,-9,-8,-53,-65,-66,-34,-8,0,-4,-19,-8,-4,3,-7,-7,-1,-4,14,21,19,26,25,3,15,15,30,26,23,29,33,19,-4,-21,-17,-63,-74,-63,-51,-13,-7,-10,-14,-14,0,-14,-5,1,0,-11,-1,3,5,-2,6,5,9,15,31,14,26,28,19,-12,-21,-16,-21,-55,-53,-72,-62,-21,-9,-1,-8,4,0,1,2,-8,-25,-16,-20,-11,-8,1,6,22,3,2,18,30,32,32,10,-10,-30,-12,-19,-51,-58,-50,-63,-42,2,4,-11,7,-2,-10,-14,-8,-15,-20,-12,-4,0,-1,10,3,23,11,14,26,37,38,13,-18,-8,-3,-12,-56,-63,-40,-57,-52,-3,0,-8,11,-2,-10,-5,-8,-7,-13,-7,4,13,17,17,22,27,18,32,27,35,29,5,-3,0,1,-2,-46,-55,-60,-52,-53,-47,3,0,15,4,-8,-3,0,13,20,18,14,26,33,40,41,18,39,28,28,28,-1,-22,-21,-9,-4,3,-30,-34,-47,-34,-49,-61,-21,6,2,0,2,0,4,3,14,13,19,31,22,36,34,28,29,40,45,17,-26,-38,-23,-17,-12,0,-38,-31,-27,-29,-55,-71,-22,-3,12,16,-4,-6,-2,1,6,13,19,27,16,30,34,38,28,31,33,14,-24,-29,-37,-22,-15,0,-36,-22,-19,-31,-56,-62,-36,-22,-5,3,-3,0,-7,2,4,8,17,27,27,26,35,25,25,25,23,8,-6,-45,-48,-31,-18,-18),(35,83,79,48,17,16,20,41,41,39,34,36,32,34,32,46,37,61,38,50,35,39,43,46,40,30,36,65,73,63,96,96,67,83,58,45,14,27,37,45,28,23,29,38,24,14,28,34,41,30,28,37,40,31,40,32,27,24,20,40,61,63,90,100,78,81,48,21,9,26,52,38,19,30,21,39,4,5,-4,8,20,15,24,25,29,28,30,24,30,46,43,32,43,57,90,88,77,73,14,22,22,40,12,8,17,1,5,18,0,-2,10,-12,13,6,5,10,11,5,20,20,29,26,27,26,33,54,63,86,78,53,27,25,30,23,28,22,-5,19,-4,-6,0,-16,-16,-1,-7,9,-4,2,18,24,13,11,20,29,38,19,18,44,49,82,85,27,10,20,22,17,18,12,3,5,6,0,-10,-6,5,-5,-9,-3,13,-9,-8,23,32,26,19,8,30,22,11,31,57,72,59,14,33,10,27,13,11,8,2,-5,-12,-20,3,-18,-15,-3,-34,-19,-20,-16,-1,12,3,23,10,28,33,4,7,28,35,55,52,18,15,21,20,10,-5,-9,-18,-16,-15,-22,-20,-8,-27,-12,-20,-8,-16,-16,-6,-4,3,3,8,21,27,15,13,30,44,64,44,7,10,13,10,6,-17,4,-20,-25,-9,-8,-20,-19,-23,-3,-20,-21,-19,-10,-9,-8,8,0,18,12,14,16,10,14,30,54,55,19,1,25,-6,8,-7,12,18,2,12,0,0,-13,-13,10,-14,-6,-28,-4,4,-5,1,11,0,15,1,6,3,6,30,46,40,19,4,12,13,-1,-3,-4,-14,0,-3,17,-5,-7,3,3,3,-13,1,5,2,-19,-9,-1,-6,8,11,22,14,16,32,53,49,43,13,5,0,-12,-10,-1,-3,-16,-12,-13,-13,-11,0,21,16,6,0,7,-19,-19,-16,-12,16,3,8,11,3,6,30,58,43,31,15,7,0,8,-1,-13,8,3,-6,0,-9,-18,-6,-23,-3,-5,4,-1,-9,-10,6,-1,10,14,7,9,6,12,34,54,32,35,18,-7,-6,1,-1,0,-6,-6,-11,-20,-13,-15,5,-19,-2,17,2,-4,-7,11,-7,-5,15,10,15,19,13,14,26,49,24,17,12,-7,-11,-5,3,2,-17,-12,-7,1,-14,-14,-13,-21,-11,-15,3,0,-5,-8,14,8,3,16,8,4,4,1,28,70,11,10,16,1,-4,-15,-5,-4,-12,6,-18,-1,-26,-3,-12,-36,-8,7,18,9,17,6,26,16,4,11,13,11,-2,9,27,36,-12,2,8,1,-9,-11,2,-7,-25,-14,4,-1,-15,1,0,0,-24,-3,-4,-2,4,7,3,-13,-8,2,0,14,17,21,24,10,-5,0,1,-10,0,-1,-17,-26,-24,-10,-9,-5,-3,-8,-15,-23,-23,-7,0,10,-7,-12,-10,-14,-4,8,-7,4,24,12,22,-5,-4,-12,-2,-6,-22,-10,-31,-37,-10,-20,-13,-10,-20,-8,-8,-30,-34,-8,-5,8,6,-5,-2,-8,6,3,16,16,7,0,16,1,-18,-12,-22,9,5,-18,-15,-24,-10,-13,-11,-4,-15,-32,-36,-26,-24,-14,-7,-21,-10,11,-13,-9,-10,-8,1,11,17,0,0,-4,-32,-23,-9,-6,-13,-3,-5,-12,-14,-19,-8,-20,-15,-22,-22,-22,-21,-19,-11,12,3,2,-14,7,-3,0,0,13,31,5,-13,-6,-48,-45,-32,-1,0,9,-7,-10,-1,-6,-12,-17,-7,-10,-10,-10,-8,1,8,12,2,-1,2,7,12,21,23,8,11,1,1,-19,-34,-36,-34,-11,-2,-3,-4,-1,1,8,10,-21,5,-11,-2,-16,5,0,2,6,-2,1,-1,12,16,5,6,13,1,-1,-37,-19,-25,-38,-43,-49,6,-6,-4,11,0,-19,2,0,-2,-7,6,1,15,-3,0,0,5,-10,3,10,5,8,14,26,-1,0,-6,-14,-28,-31,-53,-23,-4,-1,-7,-4,8,-13,10,-10,-25,-16,-3,-8,0,-5,5,3,21,-2,0,4,21,8,16,17,9,-28,-15,0,-24,-39,-30,-13,-19,14,2,-5,-3,-13,-18,-11,-9,-10,-19,-14,-15,3,8,6,-1,3,10,18,0,13,22,11,-10,-30,-1,-9,-29,-8,-28,-25,-28,8,-6,9,-12,-3,0,-10,-12,-7,-4,-28,-26,-30,6,3,24,13,9,5,18,21,24,0,4,-12,-20,-1,-12,-11,-45,-18,-37,-22,8,13,-11,-1,-2,-17,5,2,9,10,0,11,10,9,11,0,-2,16,18,14,19,5,-3,-12,-8,-10,-17,-13,-4,-42,-46,-33,24,7,-13,7,13,-10,0,3,1,11,11,21,18,5,4,21,9,14,23,26,8,23,-7,-15,-1,-6,-20,-29,-19,-23,-32,-46,-1,19,12,8,6,8,-5,9,3,12,14,6,17,0,0,21,13,3,17,29,36,11,2,-4,-7,-4,0,-19,-24,-21,-43,-58,-11,0,8,-4,-1,7,-10,-10,1,3,10,0,11,2,8,11,18,11,16,20,41,-8,0,-4,-11,-15,-20,-6,-11,-27,-48,-32,-7,-1,17,12,10,-10,3,0,-6,21,24,13,11,17,5,16,4,10,29,33,36,15,-20,-10,-7,-4),(-137,-137,-103,-44,-29,-22,7,-20,-9,1,5,32,19,30,21,6,7,32,44,25,30,34,30,7,25,8,-15,-65,-72,-85,-125,-121,-119,-87,-80,-45,-30,0,12,-8,20,17,23,37,18,37,28,6,-12,-9,20,9,0,20,42,2,42,36,0,-57,-62,-71,-114,-116,-114,-77,-34,-19,-5,11,-7,23,15,32,17,35,27,16,17,27,17,4,10,-13,9,-1,17,31,2,22,33,0,-45,-51,-61,-100,-99,-51,-28,-1,26,6,35,21,16,35,27,34,6,0,28,19,13,4,13,5,33,4,15,31,-7,38,-4,21,-17,-17,-77,-116,-63,-43,-10,14,8,17,-4,14,44,33,14,5,16,11,7,18,10,-18,-4,8,2,11,13,20,6,9,45,26,0,-20,-71,-94,-54,-10,-3,7,20,19,25,3,43,35,43,31,18,14,16,-2,0,-3,17,-28,28,35,14,-18,33,10,41,30,-19,-22,-43,-79,-62,-13,-5,1,-3,4,15,0,8,15,24,12,29,-8,16,15,13,0,4,0,5,16,0,9,6,22,48,50,3,-13,-34,-67,-51,7,-13,3,26,17,33,25,18,19,5,-7,7,7,8,-2,37,26,15,1,-13,17,6,-3,1,30,20,38,-22,0,-34,-50,-19,-12,-25,-2,22,26,0,12,0,25,15,14,19,0,14,16,33,25,3,-2,-2,2,10,6,-4,-2,10,36,11,-1,-23,-51,-34,-2,-11,5,3,5,-12,-15,1,13,6,1,-2,-5,-6,0,-1,19,15,1,9,-10,-26,-1,-13,-13,24,10,37,-10,-21,-71,-7,-5,5,13,21,-16,-17,12,-5,1,-30,-18,-4,-15,-23,0,25,4,13,31,24,3,-33,16,17,12,-4,30,30,15,-20,-36,-25,-9,-6,9,-14,17,10,-14,11,-3,-6,-5,19,12,-21,-48,-6,11,9,5,2,6,-4,2,8,10,19,44,50,5,1,-54,-11,8,-16,21,7,14,3,-1,5,0,6,-4,15,13,-13,-53,-28,18,19,-7,8,12,-15,6,-22,21,-2,11,27,24,17,-60,-35,-7,32,13,23,-16,0,-23,-33,8,-10,4,-24,-8,-23,-21,-13,6,-34,10,-20,9,-4,-1,21,-12,7,22,46,10,-31,-44,-17,1,9,18,18,-7,4,-4,-28,-9,-11,-11,-55,-9,-26,-25,-1,-9,-35,-41,-8,-16,0,-19,-10,7,-17,0,53,5,-7,-39,-10,20,-8,19,-15,-32,-6,-31,6,-23,-22,-26,-52,-24,-37,-15,-13,17,6,-23,0,-14,-3,-4,-7,15,0,44,41,31,12,-42,-4,33,17,25,18,-29,-29,8,-25,2,-22,-6,-35,13,-32,-32,-32,-22,-16,-14,-3,-27,-4,-14,-13,0,-22,-8,24,20,-14,-53,-1,28,31,39,23,10,-21,-12,-11,-12,-1,-22,-28,-21,-8,-24,-22,-9,-12,4,-19,12,8,-3,31,7,23,2,17,3,20,-32,0,6,22,43,-4,6,-1,-18,-17,5,-45,-33,-8,16,22,10,-7,3,21,22,-10,-6,0,-9,24,48,2,16,3,8,-17,-44,-3,19,7,11,16,-23,-24,4,-3,-13,-21,-19,-8,23,29,32,62,41,5,20,-49,-14,-9,9,3,6,19,-3,38,25,-1,3,-11,16,33,13,5,7,-26,-19,-6,-36,-32,-22,-5,21,46,46,61,36,40,-16,-29,-13,-14,26,25,17,10,19,28,14,7,-4,-3,-20,19,20,10,-5,15,-19,6,-27,-2,-7,6,0,2,15,24,1,7,-20,-15,-15,24,8,17,10,0,20,-1,3,-3,27,0,-19,1,53,4,-20,6,-14,3,7,-16,2,-4,-6,-13,-4,6,2,1,19,-3,-2,-14,20,30,14,26,-5,-9,11,-3,13,18,-16,23,32,34,11,-12,-25,22,-5,-21,-30,6,21,16,9,9,-1,-10,6,1,-5,23,27,-12,17,-13,23,9,4,3,-5,26,23,-5,24,47,9,1,5,9,0,8,5,8,9,4,31,11,13,7,0,4,12,28,-4,-1,24,0,-4,-25,7,10,-2,4,7,-15,16,0,6,19,-30,-1,-17,0,2,-34,-19,12,4,-16,3,10,-10,9,0,4,-5,-6,-14,8,-19,-36,-23,0,4,9,0,0,-19,33,16,-10,3,-11,12,-11,7,16,5,38,13,36,45,27,24,9,7,7,11,3,17,9,-5,-25,-14,-8,18,-21,-19,0,20,31,12,12,8,-29,7,-6,8,26,5,-15,21,-1,29,8,13,15,24,-5,15,9,20,-21,-50,-23,5,5,8,-18,-21,-11,1,16,12,14,0,-5,-19,11,-13,-5,4,2,-18,-1,9,-13,34,0,2,6,20,1,-6,-15,-44,-27,11,35,9,16,5,0,-4,-1,10,-9,-21,-7,-5,15,1,-8,12,6,23,-5,11,19,-15,8,5,-3,7,15,-14,-44,-27,4,-5,15,18,-5,-1,6,8,0,3,-8,0,-15,-7,-18,-14,6,16,22,3,11,-6,15,8,49,24,15,12,-18,-41,-51,-71,-14,0,16,15,0,25,-8,-14,-3,-1,-19,-44,-31,-17,-14,-17,0,29,20,36,22,22,32,30,21,25,-5,23,-19,-31,-24,-52,-48,-3,-21,12),(-16,14,-14,6,-20,11,0,-3,-16,20,43,8,30,-12,41,11,27,-8,43,38,52,46,27,26,12,14,-1,-18,-21,-12,11,34,-6,49,14,20,37,-23,28,10,7,25,44,39,-10,-10,28,9,-8,47,-1,6,15,26,38,25,53,45,8,-21,24,-9,-69,0,52,7,38,-39,-8,4,8,-9,-19,-6,-3,4,34,-4,-18,-9,9,-16,12,1,-36,-7,21,40,49,5,0,-23,6,2,-18,-35,20,3,17,4,52,31,8,-9,35,-4,-4,-24,0,5,37,5,43,12,-5,51,16,23,5,15,42,18,0,18,4,-27,-11,-12,28,17,6,29,7,13,5,26,3,18,-39,-27,-23,-9,24,17,14,5,16,-22,26,11,4,30,17,30,26,-14,28,10,-18,-23,-10,31,0,7,41,30,35,-3,10,-21,34,-24,26,36,2,5,12,48,35,12,34,-4,8,18,21,24,30,23,30,17,-34,4,-8,-1,-14,17,25,-21,39,7,-33,-26,-23,-18,-7,-10,-40,-4,-21,12,10,14,3,18,3,-22,17,21,19,28,3,-2,7,-21,10,18,6,-12,-20,-26,21,28,12,27,-9,2,-3,-24,9,-10,2,-5,-9,-13,2,-23,49,43,26,10,17,-16,30,3,13,-29,-14,-13,34,16,4,19,-15,-18,8,-8,-1,-27,2,-18,26,-34,-18,21,-20,-36,-4,-12,4,8,0,-7,-11,-19,-27,0,4,-45,2,-28,1,2,17,16,11,6,-5,-4,-3,-11,-19,-30,-10,-4,33,-23,-33,-19,6,-10,4,25,38,31,14,10,40,-5,10,-2,-19,19,-13,-11,10,-8,5,-31,-48,-26,1,2,38,5,-21,13,-10,4,21,-14,-23,-28,-31,8,-9,39,24,17,48,-1,-15,-17,-2,8,28,-13,4,-11,-7,-17,-2,-47,28,17,22,-17,25,15,7,19,-18,-22,48,29,14,-11,-12,13,-16,38,-5,-6,-16,-29,0,-25,-26,-2,3,-14,-44,-13,17,-21,-14,37,-23,-28,23,-29,-34,38,42,-28,-24,-2,-3,-9,10,47,-4,50,38,-26,-19,8,-29,29,26,-41,-17,0,-22,-19,-7,21,-2,4,0,-12,1,-10,11,20,13,21,-22,-18,23,-15,28,-1,3,-25,6,14,-16,-38,-10,-31,8,1,-41,-12,-1,1,1,-29,36,-9,-26,8,19,-47,-15,20,4,9,-1,-25,33,-31,-2,46,15,34,26,32,-19,-24,-8,3,-22,5,-24,-12,-25,-14,14,1,5,0,-28,-34,-37,15,0,-20,17,14,19,7,32,-31,29,-11,59,43,42,-8,-30,-68,17,-7,-35,-36,-5,-39,-46,-2,-12,15,-33,-11,-15,10,-3,-28,15,55,9,6,6,40,-4,1,18,42,36,45,8,-22,-3,-37,-7,-8,21,-4,-29,-21,-22,0,-6,-16,21,-41,3,-42,-26,9,13,9,-26,39,4,10,-1,21,-13,13,19,9,17,39,-17,0,42,-33,-9,7,-23,-19,-2,1,-18,-14,-18,0,-37,4,-21,-20,7,-4,4,37,-24,-19,-11,-13,17,16,0,27,7,7,-1,22,34,4,2,-9,3,-27,-15,-19,27,-13,-32,8,1,-28,-16,-25,-13,13,9,-8,4,-8,3,33,-15,33,-8,18,8,15,-1,-17,14,17,-28,25,-19,0,-24,-28,0,-37,-11,-1,-11,-19,-23,-2,-6,-21,21,8,26,-14,13,-9,22,9,30,25,35,-10,0,-57,-38,11,-23,0,6,-24,-3,-25,-35,-50,8,-14,4,8,2,1,-4,-6,20,10,-13,65,31,10,36,33,-17,26,-11,9,-3,-12,1,-26,10,21,-17,-29,6,5,4,7,-20,-24,-17,2,4,36,38,-9,26,5,17,15,16,22,21,1,-4,19,-8,3,-19,25,-34,3,-7,-19,-23,17,-50,-25,-15,25,-33,-24,-8,-26,30,33,33,44,5,-2,13,14,21,-3,12,2,16,-3,-53,0,-9,6,5,-22,-19,7,4,11,30,15,16,6,2,35,-12,12,2,-17,39,38,24,47,-12,30,48,-9,-11,24,-12,-10,-24,-10,-19,-31,-27,2,-39,3,10,-5,-37,14,-33,-2,18,21,-25,5,-27,22,-10,-13,3,-6,-4,25,31,-4,16,19,26,-28,-40,-9,-3,-2,-19,-7,4,-1,-25,39,32,-27,10,2,23,26,-2,-20,21,16,-5,4,11,54,6,-24,48,62,-22,-13,-25,-19,-31,-39,4,8,-36,-2,-27,-26,-2,1,-9,1,-15,-1,-6,34,0,19,1,-7,16,-2,25,-10,55,34,0,11,24,29,-9,-23,-12,-17,-22,-14,-15,-17,-4,-16,10,14,6,37,-18,3,2,-1,-18,25,22,21,-14,23,-3,-19,16,24,19,14,20,12,-35,-8,-4,39,0,-2,-4,-18,-4,-22,-55,-14,25,15,28,-34,-28,-13,37,33,2,-6,7,20,49,25,4,56,50,-11,37,0,-30,-18,-17,-13,-3,-27,1,13,-20,-26,-29,6,-7,31,21,4,44,-27,6,-8,-1,39,-3,9,29,12,26,29,-21,13,-9,4,-2,-32,6,0,-13,-12,-40,23,37,-25,-34,-23,10,-9,-22,14,-21,-19,22,-7,6,35,21,49,11,8,19,14,-16,-5,-29,-22,-13,-49,-34,14,-17,20),(40,31,16,-19,9,-3,-16,-39,-21,-17,-19,-53,-33,-48,-15,-10,-24,-32,-28,-28,-35,-20,-14,-6,-2,-22,-24,-16,-19,-62,-39,16,31,10,20,18,9,-2,-6,-38,-27,-43,-21,-39,-57,-64,-53,-17,-49,-31,-12,-41,-55,-25,-45,-27,-23,-15,-30,-26,-13,-41,-19,-15,44,-22,20,7,-25,-29,-14,-43,-25,-40,-42,-44,-46,-35,-61,-62,-28,-32,-23,-30,-48,-54,-22,-37,-20,-10,-15,-27,-24,-7,-58,-52,15,6,-21,0,-18,-5,-31,-17,-16,-46,-28,-32,-40,16,-41,-54,4,-10,-23,-8,-30,-40,-47,-22,-13,-33,-35,6,-34,-19,-40,-54,1,1,0,-4,-33,-49,-3,1,-14,-7,-41,-13,-51,-29,-2,-14,-33,-16,-32,-45,-9,-31,-14,3,-38,-15,-45,-32,-13,-6,-43,-34,-8,23,2,0,-19,-18,-31,-6,1,-29,-1,-49,1,0,-30,-20,-5,-10,-28,-19,0,-49,-21,-10,-16,-10,-14,-20,4,-12,-18,-55,15,-19,-17,-40,8,-10,-4,-9,-12,-21,-23,-5,-5,-27,-24,-7,-32,-31,6,13,-11,-25,-7,-23,-27,-9,-10,-4,-2,-18,-5,-86,-30,-11,11,10,0,-20,-43,-11,-26,-30,-4,-29,10,-20,-27,4,-2,-25,-37,-20,13,6,-15,11,-2,-27,-17,-32,17,6,3,-32,-9,-38,36,20,9,-4,-13,10,8,-39,-3,-8,-24,-27,3,-12,0,-4,-25,-14,4,-5,12,-10,17,-28,-26,0,-10,16,-13,-38,-29,-9,23,21,27,19,15,15,-18,8,17,-13,3,-28,-7,-3,12,-4,-21,6,-2,6,33,21,3,27,-6,-28,-6,-11,2,-14,-15,10,-5,46,4,8,-12,2,22,13,53,22,27,7,3,-13,11,0,-5,-7,-18,12,-2,-1,-21,28,18,-37,-12,-13,-1,-2,20,34,-14,8,12,1,9,9,24,25,11,42,6,-4,14,-12,-10,-20,-19,16,14,21,-3,-12,-10,11,-16,-17,-16,-15,-13,8,63,-11,21,30,-9,-1,22,-7,5,17,14,17,6,1,-7,-24,-40,-25,23,13,6,6,28,-23,6,12,-28,-27,-8,-15,-7,-2,40,24,29,14,-5,-15,0,60,56,20,2,-1,43,21,-5,-6,-7,-25,20,-12,-18,-15,-20,3,2,-26,-10,-25,-53,-22,7,-30,47,1,27,-26,4,32,-6,46,41,26,1,-1,20,-38,-27,-31,-19,-32,-5,-29,11,-26,-31,-15,-23,4,-10,-16,-29,-10,-4,-21,0,47,25,47,-13,-17,-27,-16,-15,28,5,5,-11,-37,-4,6,-15,-27,0,-21,-10,0,-15,-16,-5,-15,-17,-18,-24,-11,-36,-8,28,42,11,12,-28,5,7,-8,-6,-23,-35,-18,-6,-12,34,1,-9,-1,-5,-20,-19,-25,-24,-31,9,-28,-18,-14,-11,-20,-15,3,39,23,12,28,-20,10,9,8,-9,-9,-36,-22,0,-5,-10,17,-13,-25,-16,-6,-23,-13,-24,-28,-15,-44,-18,-22,12,5,14,38,31,33,44,58,15,-4,-6,-15,-30,-28,-5,-6,-12,-4,-16,3,-13,12,-23,8,-21,-4,-6,-3,-32,9,18,5,-4,-1,33,27,30,12,27,37,5,16,-20,-27,-11,-20,-15,17,20,-5,35,28,0,30,-1,-39,19,-20,-18,-13,1,8,-11,13,-25,7,30,22,60,22,42,37,9,22,25,-1,-9,13,-4,11,29,10,21,9,-21,11,-6,-17,16,13,6,-17,-2,-12,-48,-20,-1,9,17,28,24,63,21,51,49,17,12,13,-17,11,-5,12,2,-5,16,-6,12,11,13,-4,-10,-10,-13,10,20,10,-21,-6,22,25,38,16,43,67,44,27,45,19,0,6,46,38,42,-4,-24,-25,-4,18,6,8,2,4,1,38,-4,-9,11,7,-42,9,2,0,14,-8,32,38,12,17,22,39,28,16,22,8,43,-6,-13,-14,-18,-12,-20,-30,11,11,5,38,-18,0,0,6,-2,-6,34,27,28,-9,15,22,58,45,38,60,39,-12,24,35,3,29,7,-14,0,5,19,20,18,31,-3,22,7,27,-4,-30,1,6,56,30,20,2,-3,27,11,40,25,27,15,40,12,34,22,24,17,-26,-9,-33,-4,-12,-4,-8,-1,2,13,14,4,23,7,48,23,48,37,-22,17,57,22,47,23,66,57,-10,6,-10,8,10,2,9,-9,6,-33,-22,-19,-5,10,12,16,2,-20,-1,3,55,0,22,-2,-21,23,37,18,17,28,45,8,5,10,-6,13,-2,-16,21,19,0,-5,0,18,-40,-6,3,-4,6,9,8,54,45,43,-9,0,-9,20,7,36,9,9,52,63,9,-13,47,3,-4,18,14,39,-4,-50,1,-7,-7,10,-5,18,-2,-12,31,7,33,31,13,-23,-14,3,0,3,29,15,49,40,12,-11,3,2,18,10,12,-19,-36,-25,-40,-29,-3,-34,26,-7,-25,24,32,20,34,63,6,-9,9,0,26,-31,-1,7,-6,-5,-1,34,32,-7,-19,18,-15,-17,-20,-42,-25,-32,-2,-26,10,-22,-29,0,20,36,45,57,24,29,-23,-16,-4,-10,-8,-26,-10,-16,-12,0,0,41,-4,-5,10,-25,5,0,2,-18,14,27,-9,-19,-22,-26,28,44,49,23,8,29,-21),(9,70,106,54,19,31,15,3,-51,-16,-36,-41,7,13,2,-44,-34,-4,35,-45,0,-62,-53,11,-10,2,42,27,62,48,-3,-18,60,106,25,62,-30,8,55,-34,-1,-13,-42,-52,-67,-53,-63,-60,-4,-31,-10,-26,-8,9,-40,-22,-4,3,73,51,-22,15,-1,20,105,90,26,13,58,5,-45,-48,-29,-7,-73,-6,-13,29,9,-6,22,17,-47,24,28,2,0,-10,-15,-9,-11,0,22,-19,48,-5,63,83,58,46,1,13,18,5,-52,-50,3,34,-25,-37,14,5,11,-32,32,47,3,-17,45,43,3,-16,-34,14,53,-11,46,-18,92,36,-12,41,30,-54,-31,-64,26,-79,18,-15,-51,28,-34,-12,24,-24,29,9,36,22,20,16,24,38,-17,22,41,-17,48,21,92,-13,27,-8,-48,-24,-59,-79,-7,-46,2,-16,3,4,33,-2,0,-27,-21,0,10,63,38,-35,-30,5,15,-8,-40,29,-13,8,65,9,14,5,28,-14,-37,-24,-68,-51,-57,37,-44,-46,14,-12,-39,-46,-22,-17,-3,8,-22,24,30,30,38,23,71,-23,15,20,-8,32,9,-35,-50,-22,6,-24,-45,18,46,0,0,31,23,20,58,27,-10,-3,11,55,46,-28,21,-7,27,26,2,-20,52,39,77,51,45,54,-41,-15,-13,-34,-3,-23,-42,18,-38,-41,-11,26,3,25,1,39,25,11,9,-15,-43,-18,-23,-11,16,8,59,-18,60,-9,56,-39,-22,-10,-20,1,-46,4,25,16,-21,-63,-1,-25,-44,-2,-36,-56,-46,32,-47,8,-22,2,13,-25,61,37,0,-32,33,78,73,14,7,12,40,-19,56,-18,9,4,-3,20,10,47,-14,-44,-36,-16,-30,22,-36,-4,45,47,27,27,44,2,-35,11,56,11,31,-11,34,42,47,41,38,-15,-27,65,31,36,-44,4,60,-57,-49,6,5,54,54,-4,-21,-19,-18,-21,66,-10,-17,31,65,-19,21,26,-33,6,-20,48,51,42,-13,30,-15,33,36,-21,-12,-20,39,2,-24,9,-36,18,12,8,-41,-43,-19,-24,5,-6,32,0,33,-24,-25,-57,-15,-8,23,0,17,-40,-49,53,-9,6,5,29,-16,63,-26,-3,-4,47,-2,-49,-46,47,-25,-19,9,-6,18,47,62,38,-39,50,-34,32,-21,-46,-51,7,-35,-21,-29,45,68,-40,-35,-23,-3,-23,9,13,-45,14,-29,36,70,-53,26,-50,58,-14,-39,-30,-21,-20,51,-36,-12,-20,-2,2,-12,-6,-21,46,-55,25,-7,-17,-37,25,-9,-18,73,-1,52,15,68,-5,0,-31,-25,-52,-19,-48,-50,-45,0,72,-49,4,-25,18,-35,-31,22,-37,-8,-17,33,64,2,-48,-11,25,56,29,-35,-6,-15,-32,-37,-61,-40,-66,-8,34,-32,-5,39,-5,31,-2,-4,44,-28,49,50,83,59,-21,39,28,48,49,26,-20,19,-25,16,-48,45,24,-80,-28,63,25,30,37,-5,-5,-36,-16,-46,49,46,63,-16,-26,24,29,19,-26,32,-32,40,62,-32,34,-27,60,54,15,-15,-46,-51,-4,55,19,-39,13,-27,-9,18,18,-3,-34,51,-29,-9,10,-46,2,-29,-43,-20,42,-24,2,-18,24,37,-59,-14,7,-17,-1,-24,-16,24,0,-36,-11,14,49,-20,23,-31,-29,43,6,-32,-35,13,-14,-25,-17,-31,12,42,32,-3,50,-11,-54,-14,32,-46,-55,-2,10,22,-35,-59,-22,6,36,-24,-11,56,-61,11,-45,-36,-28,-34,-43,10,-7,-45,-64,15,25,10,0,-26,-19,30,-5,-52,-89,-51,-19,70,-19,-59,15,-48,-9,0,14,8,-3,-19,-52,-46,30,1,19,-14,-2,28,38,-8,35,-27,26,32,30,-65,-62,-30,-27,6,-43,-12,-18,-61,-29,-68,-40,8,-25,29,11,17,7,-7,-3,-24,-9,15,-4,41,-11,50,-3,9,41,-50,0,-33,-33,-35,-74,-53,11,86,-2,36,-71,-13,-8,-25,-13,5,-65,-19,29,33,-54,-11,-17,-28,13,3,54,-24,49,1,-4,-4,-61,-1,-92,-69,10,-42,43,-18,34,-30,3,-17,-38,-22,15,-66,18,-29,17,-13,-39,-16,-23,49,6,30,-20,-6,12,-54,-45,-17,23,6,-30,-75,19,51,-34,0,0,2,-21,11,-7,-20,2,-13,2,-2,-43,-51,-43,-23,25,-10,15,-24,-20,-18,-14,4,-46,-23,-2,-13,-7,-50,-18,13,10,-11,61,45,-40,-36,-68,-26,4,-63,10,4,-61,16,-1,-26,-24,11,-42,-33,-68,6,-56,-38,-38,-23,-3,-45,-58,7,17,-16,31,57,-38,44,30,-36,-22,-23,12,-31,-29,4,29,-39,11,-24,27,5,-31,22,19,-28,-14,37,-36,23,-3,-32,-35,40,63,47,52,42,-4,58,28,-37,44,-31,-49,-21,16,22,-10,-16,-42,-19,-31,24,23,34,2,-6,-59,-48,31,-31,-10,12,1,66,67,0,36,-22,33,68,77,-5,11,44,23,-18,16,-19,-37,-34,-50,10,-54,-6,-59,-25,-1,13,-53,-49,-5,6,-39,1,2,66,13,35,65,32,55,25,47,19,80,31,10,5,-39,-26,-26,-38,29,-56,-2,0,-11,-28,0,49,17,-2,-9,-67,-18,16,77,68,7,31,10),(71,99,54,43,38,-4,16,21,7,4,-35,-43,-40,-42,-17,-54,-32,-63,13,22,-25,-1,-18,-25,7,14,36,-3,47,51,68,76,42,118,44,-13,43,-44,0,1,-9,-14,-38,-42,-74,-40,-67,-23,-49,-11,9,-44,-63,19,-22,-6,-27,20,14,11,53,37,61,85,98,71,14,3,-25,-33,14,-8,-50,-61,-11,-83,-25,-72,-22,6,7,-17,31,-26,7,-8,-5,-46,-38,3,-46,3,48,46,50,43,48,-8,18,-11,-5,-49,19,-32,-38,1,-29,-50,-8,-26,29,3,-34,-38,-16,14,-3,-20,-2,-31,-49,-4,-3,31,-7,37,54,66,85,14,27,-10,15,11,-31,6,-3,-17,-35,-40,-10,-54,6,0,-25,-50,-14,-2,20,-37,-49,-25,-12,-28,-13,-8,-3,22,68,11,3,-4,-1,-2,48,43,17,0,-15,-12,2,-51,-28,-9,-39,-54,-24,-46,-38,-13,0,-13,-30,2,27,10,-31,32,-24,24,19,77,30,22,-18,-25,11,36,16,-51,9,-33,19,1,-18,-15,0,-48,19,-48,-48,-23,-44,-10,14,-36,-31,-41,-2,-2,-26,12,72,21,30,18,1,35,24,1,34,38,21,-50,-60,-14,8,-32,4,-38,-9,0,18,-9,-22,15,13,12,1,-13,-2,-3,-38,2,-17,-7,20,8,1,2,9,-2,-12,-26,-49,-10,-27,-38,8,-16,-20,-37,-18,12,-23,15,-36,-56,14,12,-16,-15,-31,-22,-34,11,26,26,12,11,25,9,15,-44,20,-22,0,51,24,19,-19,28,-22,-5,-26,-30,-9,24,16,-52,4,-31,9,-4,-30,-60,13,-33,-15,18,-3,9,-14,2,10,18,55,43,35,41,-16,22,-20,-45,-4,-5,-6,-34,-33,56,44,0,-25,-20,-6,-33,-41,-11,-43,-23,1,48,60,15,32,56,4,21,17,-2,15,29,26,20,2,11,35,-32,-31,-53,1,23,35,19,13,6,-5,1,-17,-52,-89,-3,9,61,14,-20,-24,57,18,-15,28,-37,25,16,-26,-5,-7,9,13,-57,-14,-25,-10,18,20,54,-5,-16,-26,-26,15,-6,-83,-39,72,44,35,-2,40,2,-5,34,6,26,2,52,30,34,-17,29,17,-56,-24,-7,-28,-5,-8,-4,-25,-47,-11,21,1,-9,-8,-32,-6,53,68,56,37,10,39,1,26,5,5,-12,54,-1,12,7,4,-32,-26,-10,-32,-6,4,0,37,15,3,5,-32,16,-63,0,12,44,18,42,2,52,7,-17,25,-18,54,13,-1,20,-40,-7,-29,14,12,-16,-27,-1,-31,-29,1,-54,9,-35,-19,-30,-21,46,-3,69,35,-4,-14,43,0,36,24,1,5,-4,-39,25,-19,-5,14,5,-36,-23,-22,4,-16,5,-3,5,-63,10,-27,-50,-19,-8,46,49,41,12,57,8,-14,4,25,40,-2,20,5,-5,-19,-50,14,-34,-7,-8,-41,3,-28,2,-25,-16,9,-28,-51,-4,-49,0,1,37,28,26,-2,41,12,44,0,23,-43,-8,-9,7,-20,28,-6,14,-12,-7,-7,-18,-12,-30,-51,-33,-22,-20,-13,-6,-8,-6,23,70,41,41,74,0,49,-6,-2,6,5,13,-7,23,-12,2,-47,14,21,14,-33,-14,23,-32,-35,-36,3,22,-39,-34,28,14,38,72,-9,15,35,5,17,36,-36,3,37,-42,1,27,-4,-2,15,22,-2,-29,-11,-34,0,7,3,-31,-9,-12,-2,-10,2,-9,88,-5,30,19,9,21,7,22,5,6,-16,-19,41,3,46,41,38,19,-28,0,-2,40,-15,-42,32,-38,2,-42,-10,13,17,40,38,0,0,-45,34,43,30,20,-11,21,54,-9,0,1,29,37,38,32,58,45,16,14,14,-55,28,-5,-3,17,24,31,36,33,48,55,5,27,16,-8,21,28,-33,37,51,-2,-18,10,0,25,59,63,10,-12,2,12,18,-1,11,-25,-7,-27,-20,-6,58,2,-9,21,19,32,-40,11,47,36,3,10,-8,35,22,-1,5,18,-19,-6,1,-21,6,0,1,-3,6,-13,-2,-15,39,41,57,7,48,2,19,19,2,2,21,5,23,41,32,-29,10,38,-3,-13,-5,-25,-15,15,-4,-9,26,-5,18,-15,-45,-60,-20,50,10,-8,-2,-1,2,-18,25,-18,-32,24,55,24,12,39,44,40,-22,-24,-12,-55,-8,-16,-9,21,0,10,31,26,3,-11,29,84,0,25,11,10,-4,16,12,25,-4,15,22,35,39,-1,27,8,1,12,14,-11,2,-30,-18,-6,-11,18,-22,-20,-15,-1,48,54,37,-47,-16,-10,-30,21,-47,-16,-22,-51,-19,0,34,-10,22,16,40,-12,13,-1,56,41,-1,19,-14,4,-5,3,-15,19,37,39,17,-21,5,-42,-9,52,-9,4,-36,-36,-18,32,6,24,-3,-6,4,-19,9,24,-39,-52,-1,0,-19,6,-41,-21,23,71,62,49,-7,-18,-39,-3,-16,-21,-40,-51,-42,-33,-66,20,44,55,-14,31,-12,-19,-44,-29,-53,-29,1,-9,2,-37,-34,22,-21,37,25,29,29,4,24,-29,4,18,-65,-53,-44,-91,-23,18,41,17,1,42,-3,32,29,11,5,4,8,5,-15,2,-14,24,15,20,54,39,11,35,9,26),(61,57,40,9,-13,7,-28,-28,-44,-25,-29,-50,-28,-4,-26,-41,-34,-42,-35,-60,-31,-48,-45,-19,-52,-10,-18,-12,-41,-2,15,8,96,77,28,6,-43,-43,-42,-33,-47,-32,-43,-50,-29,-20,-38,-33,-8,-20,-57,-7,9,-19,0,-32,-39,-36,-16,0,-15,-16,-22,14,59,78,6,-22,-19,-52,-54,-20,-59,-25,-50,-28,-18,-34,-5,-5,-40,-23,-53,-32,-22,-14,-26,-9,-8,-36,-18,8,0,-26,-9,14,61,57,6,-24,-19,-47,-29,-51,-35,-38,-55,-45,-23,-53,-25,-2,-38,-14,-27,-23,-18,-11,4,-7,-13,-5,-18,-35,-6,-40,-23,-19,51,9,-31,-10,-21,-18,-27,-60,-34,-37,-31,-47,-11,-29,-56,-14,2,-11,0,9,-2,-15,-14,-18,1,-31,-7,-17,1,-18,-31,-34,90,-3,-14,-23,-51,-41,-34,-41,-50,-6,-60,-23,-34,-35,7,-17,-27,17,12,-27,-35,-2,3,-18,-21,-50,-23,0,-13,-14,-16,-6,33,20,10,8,-31,-60,-36,-15,-48,-19,-51,-52,-31,-12,-30,-19,-23,3,-36,-39,-4,-16,-35,13,8,2,-14,-19,-22,8,-32,-17,31,4,-6,-25,-50,-24,2,-27,-17,8,-54,-29,-46,-4,-2,-27,-25,-18,-19,-20,-34,-22,-3,-22,-16,-37,-8,1,-25,-25,-7,2,2,9,-33,-26,-42,-33,-29,-28,-34,-19,-43,-16,-15,0,-19,-26,-18,-12,-4,-18,-8,-10,-15,-17,-34,-10,-3,-29,-17,-13,-27,-32,60,-21,-27,-19,-49,-4,-51,-13,4,16,-5,9,-31,-24,-11,14,-11,0,-20,-31,9,-21,-28,-11,2,-25,-19,-34,-33,-27,-10,-43,52,-20,-19,-39,0,-25,-10,-11,-3,22,10,14,2,31,17,18,-18,-20,5,6,30,3,10,12,13,-20,-25,3,4,-9,-33,-7,33,-17,-5,-19,-12,7,18,18,10,-15,-2,-15,27,21,-7,10,-2,13,8,17,36,17,16,8,2,-34,-46,-32,-5,-23,-21,-5,23,34,-31,-29,-20,20,-3,23,-28,0,-10,-9,22,23,2,-6,-7,23,38,2,22,-20,-13,19,9,-12,1,5,-5,0,-27,16,36,-5,-18,-21,-11,17,0,-23,-22,17,20,19,7,-22,11,14,-6,9,-8,10,12,10,24,-7,-23,-11,-11,5,-22,-12,-35,8,10,27,-20,10,-18,-8,23,-22,-4,-6,0,0,-11,18,13,5,-7,12,0,0,0,5,3,11,13,-15,-16,-30,-16,-8,-11,11,56,-6,-1,-32,6,1,-11,4,4,-15,12,-3,0,18,8,10,-12,-27,7,2,-13,-15,17,8,-34,-25,-7,9,0,-19,7,5,52,25,25,-32,23,-13,-14,-9,-5,-2,15,-26,0,-15,-15,21,-8,-10,-31,1,-10,0,-19,-8,-33,-12,-9,8,-20,-16,1,57,52,46,22,-2,20,-15,-13,-15,-23,-23,8,-32,10,38,28,16,-5,-13,7,-3,1,-1,-28,-3,-7,5,8,-10,-18,-13,-3,19,79,51,3,0,-30,-3,7,-2,20,32,-7,-5,4,3,13,1,-19,-31,-24,-10,3,-7,-1,-1,13,-21,-22,-20,-2,25,40,54,56,80,41,7,4,-5,11,14,-12,-16,-14,-20,-9,17,-27,-19,-3,-31,8,11,-16,17,8,-1,-22,-27,8,-1,5,11,38,38,29,98,18,36,-2,-19,-9,-14,-11,-19,8,18,-24,-21,8,-3,-4,-29,31,15,-11,0,-12,-1,-1,0,18,4,41,27,52,30,47,67,26,12,11,-9,-11,15,23,-4,0,-10,-2,3,-31,4,5,4,-4,10,18,27,9,-9,10,11,6,25,24,32,20,38,21,31,61,24,10,-2,24,28,-21,-26,-15,-2,-4,16,26,-26,4,-18,14,-1,6,-21,-11,17,-11,-21,10,3,21,35,15,5,4,35,79,25,66,19,-8,-2,-9,11,-18,11,5,-17,-12,4,26,27,-15,-1,11,-13,14,15,17,-15,0,43,2,19,36,15,7,-3,28,71,21,-9,-24,31,12,-5,9,-7,-8,13,-10,-7,-6,2,-13,-19,18,8,24,-28,-15,7,-8,30,40,22,11,21,25,18,61,84,78,32,3,-34,20,-21,-14,-9,-19,25,5,12,-35,-26,2,28,-10,2,0,0,-24,-8,32,16,32,-10,14,-3,-27,-7,4,42,73,28,-3,8,-1,-2,-1,4,0,-5,11,-31,12,-13,10,18,-4,-10,2,-5,-2,3,40,31,46,-7,-6,-1,0,-4,-9,23,46,33,42,15,-3,6,1,4,9,5,-10,-15,11,20,-1,26,15,-3,-30,17,-23,2,8,16,-4,33,-8,1,13,14,-7,-8,53,46,21,42,8,-17,20,-5,-29,17,-17,24,15,2,2,-9,8,7,-6,-25,6,3,45,28,12,-2,9,2,1,5,-14,0,42,54,44,29,18,-4,21,7,11,7,24,13,7,37,22,-5,-3,-14,2,13,-15,42,56,3,0,-13,-2,-3,25,-31,14,-5,-10,37,89,43,-10,-5,9,13,-16,9,13,19,21,25,7,-14,6,-4,12,6,-14,38,47,18,-31,-23,-35,-2,-9,-31,-14,-29,3,25,30,38,-7,30,-41,-13,1,-21,-14,-38,-3,11,7,-28,-24,-11,-6,-7,9,8,6,-1,-10,-23,-32,-3),(0,-11,-36,9,3,9,20,-62,-4,8,-43,54,46,59,-34,12,64,8,23,-55,30,14,-4,0,26,-15,-7,25,8,28,-30,-29,70,1,-49,3,-45,-2,-14,-21,-29,-7,14,64,16,17,-34,-69,13,-25,-37,-25,-11,-23,38,-21,-24,-37,9,32,26,-5,-72,-7,-6,19,57,46,-12,-19,-13,-8,-11,30,30,0,-4,-30,54,-24,-25,41,-50,-60,17,36,-38,46,31,-2,-2,-30,39,0,-34,-39,22,25,-4,-4,22,-42,-4,55,13,-41,-36,-17,0,-25,-27,-12,10,-29,-16,-54,0,-36,-83,45,7,-47,-64,23,38,-32,57,-22,16,24,1,-10,36,-32,-55,-42,-19,-1,28,-3,-18,2,-6,-8,42,36,-26,5,-41,69,22,-27,-53,-19,8,52,26,-22,36,17,70,32,19,-63,-36,-18,-15,-48,-23,18,6,26,-16,-2,-20,14,-49,-46,-32,31,-30,20,-33,-32,-18,-50,-77,0,-72,55,-24,11,-17,-15,-17,0,-37,15,-3,14,11,-24,-13,-14,2,-27,-23,5,-18,4,11,-49,-14,-7,-67,-28,-18,-19,-63,-26,5,41,-48,32,-43,-56,-53,-31,-36,13,-61,-39,32,-9,-17,-40,-65,-4,3,31,0,-19,-35,-40,3,0,-34,-47,44,-2,-53,-5,-11,7,6,1,28,33,16,-59,11,-3,-40,-55,-6,21,-4,-33,-8,-53,6,11,-21,3,-17,4,-2,-8,-11,-61,13,-24,-18,-12,10,-13,40,-39,-24,6,32,-14,-68,-2,15,4,32,-36,-33,-31,35,1,-1,-42,57,-16,-11,-20,-45,42,-1,-30,24,14,13,14,40,-25,17,-18,41,-38,-52,-49,13,-40,12,-29,39,-48,26,10,-50,40,5,28,23,-56,55,-25,-53,36,27,51,43,33,25,-32,36,7,-11,-5,1,-30,-37,23,-47,-27,-6,13,51,7,1,33,-19,85,-27,44,-9,18,28,-26,-20,5,-15,-27,-19,14,21,-3,-9,-53,-12,-32,15,1,5,1,-5,30,-8,34,-42,-2,-84,25,-7,-32,64,-18,-22,-23,21,40,22,0,-4,13,58,-4,-47,-56,47,-80,-9,-26,-17,53,25,-67,14,-39,9,17,-5,-11,25,22,13,0,29,-25,-6,-22,-34,-26,17,-25,-9,-41,-4,-32,-9,-18,0,42,-13,17,85,-29,35,-11,-19,11,6,7,-16,17,44,-10,-5,-26,-14,13,-1,-7,-19,15,5,-36,7,-15,24,14,15,-2,23,13,-43,-43,76,24,-40,-45,-15,28,-24,-23,13,-6,66,-36,49,27,36,-1,-10,-10,-10,-11,20,-24,42,-27,-48,-29,51,-44,-28,19,-20,-1,-22,-6,1,-31,-4,-2,-6,5,-2,-18,-14,-32,3,35,-33,-37,-49,-44,-17,-3,-26,-39,24,42,-23,-18,22,-1,44,0,-37,-52,81,-35,13,-67,-12,33,9,-6,23,-9,-31,19,12,9,-38,-41,36,-56,61,-50,51,17,-24,-7,-25,18,60,70,-30,11,-3,17,9,56,0,-34,37,32,24,0,-54,12,-15,-52,-72,33,-10,-36,-28,-17,-43,-4,3,53,-44,-3,16,40,-21,-7,-43,-8,74,25,33,53,7,-4,-43,-62,23,-42,15,-56,27,-41,-9,-90,-33,-15,-37,-34,54,-22,-8,-18,35,21,-5,-36,-11,-30,13,71,35,6,-30,-16,66,49,-15,24,-53,-36,-31,23,-26,12,22,55,24,-15,-17,48,35,73,40,-9,0,-16,-46,16,20,0,31,52,-36,16,7,15,7,22,-20,0,-5,0,-35,-28,-10,-13,-36,53,55,-19,48,-29,-21,-25,39,12,3,29,-60,2,-16,-14,-29,54,13,-13,32,27,-21,22,45,-22,-46,-20,-14,12,6,34,60,17,41,-7,-18,16,26,44,-25,52,-6,43,19,15,39,-19,63,33,39,-5,-33,-23,13,1,28,-1,56,35,-48,-22,-38,33,-2,37,21,-61,0,-14,-37,-29,-28,35,53,6,29,8,3,59,13,12,-8,32,-28,-48,63,10,65,36,4,40,30,-9,-5,11,-44,52,0,7,-49,-16,-35,43,28,46,16,3,51,76,-25,58,16,13,25,24,-7,20,36,16,74,-15,43,26,-41,51,-5,-17,-33,-9,-45,-30,-24,-5,-41,-18,27,43,28,-34,37,35,43,41,23,58,7,34,33,51,28,-2,-4,24,2,26,27,-17,-10,-26,-41,-62,-15,-13,-31,35,-26,-17,-37,60,41,4,29,10,-17,10,2,36,-53,7,24,0,55,10,22,24,15,-1,-32,46,24,-11,16,-50,12,-22,-18,-27,32,-32,61,-32,36,33,67,15,56,-15,-5,28,61,-11,-66,7,47,9,83,65,93,50,7,-14,28,-6,-22,45,-12,36,4,26,-12,-37,-23,-2,-35,2,-20,-39,27,28,58,-33,-49,39,58,26,-42,-12,-27,62,6,-4,46,-1,-25,62,40,-25,10,8,-37,7,-10,-6,-16,9,-7,65,1,-16,-40,-20,1,43,-26,6,30,-45,-34,-27,-33,-29,31,51,-35,-17,36,33,7,-34,-2,-5,-34,20,0,44,-31,-37,-13,8,-1,62,-5,-60,3,-31,-57,58,9,-34,52,7,-57,38,17,-11,36,-1,4,30,-1,22,-22,0,-47,-24,-11,-5,1,-1,49,-36,51,-30,-63,-53,-47,-91,-24,-3),(-41,-15,-34,9,-14,-7,25,14,12,5,-4,0,53,-21,19,-29,-38,-49,43,-21,-5,9,14,2,33,44,39,22,-37,20,-49,7,-36,0,-46,19,-8,5,22,22,-38,45,46,-2,2,-1,-45,-32,45,60,52,37,11,51,11,44,11,24,-13,-34,-24,9,27,-8,-72,-64,-10,2,18,-35,-43,48,23,29,7,31,49,21,-7,-9,-26,37,37,-6,8,8,-33,-21,18,-36,13,15,-20,-27,-24,-37,-70,-73,-15,7,-2,29,7,13,47,27,14,0,3,7,60,0,22,0,12,4,-22,6,-40,45,5,-1,0,-9,-42,-59,-12,-35,7,-60,-10,-10,-28,10,5,32,24,9,-15,28,1,-10,23,-32,36,25,29,27,22,-27,-1,25,-9,0,28,38,1,14,-29,-47,-7,-65,14,-22,6,14,36,0,5,4,34,-18,41,-23,18,-23,-1,-6,47,33,49,-22,-4,1,34,25,11,50,-38,-29,-29,37,7,18,-44,-51,25,15,31,23,17,39,-17,-32,-19,30,42,27,10,22,36,17,-29,12,25,14,7,26,15,8,-29,-29,23,2,-25,-38,-24,-38,-57,-33,-37,42,31,25,7,27,36,47,0,-24,38,21,30,4,35,34,47,-20,2,-18,44,16,21,6,15,-11,13,25,-55,-28,22,-25,-33,38,63,12,13,60,47,57,41,14,15,-29,27,-18,-3,-49,-13,-30,31,-3,43,6,6,19,-14,-38,8,-33,-40,-3,-27,-46,16,-7,-53,26,-6,49,1,-23,-30,-38,-28,-5,-19,-43,19,-51,4,11,16,0,0,-4,22,3,-4,-8,12,-23,-54,9,-3,-15,-5,11,-58,-63,-12,-39,0,4,-11,1,25,16,-14,30,16,-9,7,14,19,24,41,27,63,6,1,26,11,12,-34,33,29,-27,-57,11,-7,-46,-36,-22,-44,10,6,-4,50,-40,-4,-12,-11,3,18,10,14,6,-26,5,-24,15,-14,-2,11,-5,-10,12,1,1,-46,-26,-26,26,-66,34,-61,-9,-25,21,37,7,-15,15,29,47,15,-9,-20,-29,1,29,-8,-4,24,-28,2,6,-22,1,19,7,-57,-45,-40,17,11,27,-26,-38,-10,-13,46,10,54,-12,23,6,34,-46,9,12,-9,39,43,46,4,-40,38,-6,-19,-63,-14,-3,0,-2,-24,-18,4,-2,-22,-66,32,-30,-2,-15,13,0,-16,-32,9,26,5,47,36,34,-16,12,-6,-62,0,5,2,-24,-2,-38,-19,-5,-37,3,-51,-7,35,12,6,9,13,-37,39,63,-4,14,43,-1,2,24,-13,-8,11,41,1,9,5,-6,4,-65,2,16,-31,-35,-15,-26,-11,-7,-6,29,12,-38,36,30,0,-19,25,84,63,74,44,42,63,15,-12,-26,59,-4,10,-25,11,4,-15,-2,-4,-14,39,-39,22,-31,29,-13,-52,-25,33,4,-13,-24,23,28,-24,38,16,8,4,58,46,-18,-72,-8,8,23,-30,-8,-31,-41,6,46,-48,5,40,20,-3,-35,-30,-17,-11,4,-36,31,20,24,-4,54,61,-5,53,-13,14,43,-30,-18,4,-12,21,-40,6,9,-10,8,-2,-37,17,30,12,-41,-10,-15,-3,3,-10,-37,11,-41,28,-4,87,43,-39,-56,12,12,-64,-19,47,-15,-56,-25,-31,-12,11,-31,65,-10,49,3,3,-43,-18,-24,-2,1,-28,9,21,-16,54,-13,17,-19,26,0,-10,4,26,-7,11,-28,4,28,-53,-16,-17,-26,5,-22,-48,-15,30,-14,-2,47,29,4,23,-32,17,21,-14,13,5,4,0,-23,29,-33,-31,10,27,-12,45,-10,-38,1,-34,13,-35,0,-39,-26,-5,13,-11,4,-27,-19,12,32,71,6,9,-19,1,-4,12,3,-54,-50,-4,-26,9,28,-24,3,-21,-34,-43,-46,22,-13,-21,45,-25,-7,-7,37,4,24,18,33,42,-23,20,2,65,-26,10,5,-31,-29,28,20,17,3,-8,32,25,-25,-2,-40,-34,12,14,6,-44,-49,-28,-17,32,-1,19,39,32,-24,22,-21,-9,-19,31,-18,-11,-53,-4,3,-1,60,12,-9,24,-56,-40,16,-20,-51,-35,-20,-35,-34,-50,-39,2,5,17,27,-55,-7,2,-26,7,21,-25,6,-88,-40,-6,-29,-13,8,5,19,-30,-34,-13,-27,-5,-1,-23,30,-33,4,17,-5,24,-21,-12,45,27,25,35,-27,20,27,-51,-27,-43,-24,-1,-29,-21,16,-3,1,-42,-13,-54,-21,-9,-54,30,-21,-24,11,14,-10,17,-11,26,19,-1,-55,-46,-24,34,-6,-36,-105,-70,-9,55,-10,-15,25,-14,11,17,5,-21,-67,28,18,12,29,-10,7,-40,-2,2,27,-16,-15,-17,28,-1,42,-24,8,-43,-9,-8,-32,-8,16,-2,18,-10,-12,44,8,0,-20,-45,-3,-20,7,12,8,27,26,-45,13,50,8,-22,46,2,-13,-3,-35,-68,-54,-2,-6,-19,-18,32,20,22,42,11,23,-21,29,26,-25,-11,-8,20,5,2,-6,-5,14,-21,-15,26,2,29,-25,-65,-56,-68,-27,-38,-25,44,-23,-17,4,-8,62,20,25,22,-5,-62,13,5,-10,7,19,-30,22,-11,43,15,-45,23,-3,-26,-14,-1,-89,-26,-73,-2,-39,-24,-21),(133,71,58,-6,-51,4,-42,-40,21,-30,16,-19,-4,-57,-43,-15,-14,25,-26,49,-28,30,-4,-10,-19,-26,20,-8,3,8,29,46,52,71,52,17,31,9,3,29,-17,-42,0,-25,-5,-69,-1,-11,-35,0,22,-14,28,-54,-39,35,26,19,-21,-23,-38,-18,22,0,97,20,-12,-1,-19,-45,1,21,-49,-5,16,0,-39,-51,-54,8,-11,23,52,8,-42,2,9,26,55,-52,19,17,-16,-63,24,1,73,37,26,7,-22,23,0,4,-14,-67,-29,3,5,-25,-3,-3,-25,-17,47,12,24,22,-30,-31,-16,-7,-3,7,-19,8,-60,28,87,49,25,-41,-32,35,8,-46,-44,1,-29,13,29,27,38,-14,-52,-10,-8,-13,-32,-13,-1,-18,25,-25,-5,54,-32,-26,-61,-15,23,66,0,-16,16,-69,8,15,-21,-36,-3,13,-21,21,20,9,-22,0,34,18,73,-18,4,2,42,-5,42,10,-8,-4,20,-24,102,28,23,-31,-81,3,-16,-26,4,-27,0,-2,21,12,13,36,-30,-2,-5,20,-19,-18,-13,45,20,16,5,-23,11,-34,-48,18,-2,-45,-28,-39,-2,-12,-15,6,9,-51,-15,6,6,-31,-52,-1,-26,-49,10,35,38,-27,-49,1,-34,15,9,21,-19,-10,-2,-23,-24,-2,0,-70,-35,59,-7,-9,-37,-16,-29,-34,-48,-21,-36,27,56,0,-22,-35,-2,30,-17,-49,16,20,-44,-9,45,-51,-16,-12,13,-28,-63,-63,-27,0,6,-3,-20,-23,-62,24,-5,-7,32,26,19,-52,-14,-5,-42,-19,0,-11,-8,-39,49,15,17,38,-3,-13,71,4,25,7,-14,-3,-30,-10,18,47,21,-3,-19,-66,-8,-56,-53,-3,53,-6,-38,37,-30,1,-16,11,18,-17,-4,36,15,-39,69,43,-65,-75,6,-70,-11,5,-11,11,42,-16,4,-16,26,-32,-55,-15,37,-33,-20,38,9,2,28,-1,3,-29,-2,-32,54,11,102,10,-25,-67,-55,7,-35,12,28,5,22,-12,3,-17,38,-17,-39,18,-9,-37,-52,-43,55,-27,8,63,21,34,-32,5,-38,21,63,56,-7,19,8,35,10,0,25,33,-14,37,2,-30,-23,55,4,30,32,43,50,-44,3,21,-14,28,-4,-8,-17,6,39,-27,14,18,-14,-6,-11,8,-54,40,-43,36,-49,-29,23,-11,48,-28,13,9,52,12,-21,-6,-6,-44,-10,17,-9,7,0,-6,-41,8,-19,-36,-11,-34,-19,26,18,12,0,-14,-27,-12,-24,-6,39,-20,-24,53,17,-40,6,-1,15,19,-18,68,-14,57,-7,8,18,-7,2,28,-3,-87,-44,-60,-21,0,-8,33,8,-27,35,32,11,24,0,30,13,22,61,28,-25,-45,-1,9,-46,16,-41,2,36,-34,70,62,10,-7,-10,-32,-50,34,15,-8,-25,9,-8,-44,-20,-17,-27,-14,58,40,49,-29,20,20,25,-22,8,-11,62,-38,11,-32,21,34,-12,-39,-3,-64,-9,-35,-12,-22,-40,-22,25,-14,2,-9,-68,-21,23,36,45,-29,13,11,3,31,-46,-25,-51,-12,-2,-31,43,24,-15,9,-24,20,-20,-21,5,49,-13,-26,9,-13,16,-53,11,-47,37,20,-8,6,58,49,-31,57,34,16,9,44,-27,-19,23,19,-6,17,31,-21,2,-25,-15,35,-37,-56,15,32,-63,-37,24,-36,-34,8,-17,47,12,56,42,-31,30,-21,-13,-9,-10,10,-6,10,61,-9,25,-17,-26,-83,-24,41,14,3,-22,-32,-65,-36,8,-17,56,-16,-22,-5,21,-23,-28,31,30,36,51,18,-17,-12,-73,49,35,44,-41,-43,38,-57,-31,-18,-41,67,-26,15,-33,16,-23,-12,51,-23,52,9,-32,15,0,-58,51,1,18,-31,-31,6,-1,-19,44,3,-18,-9,-19,-59,6,49,25,-21,42,0,18,45,12,29,23,-10,8,4,-27,13,32,39,23,-31,-10,1,19,-39,-24,21,80,17,40,24,-2,16,-3,18,-29,4,-32,11,33,5,-21,39,55,12,-40,-55,-28,39,2,52,14,74,11,-28,22,-6,-77,8,-52,35,6,42,-7,-55,0,-12,29,-43,14,-40,-31,-19,18,9,16,-42,-3,35,19,44,6,-29,-30,33,7,45,-27,-6,37,-26,-11,4,96,36,28,-8,-34,16,-37,-14,29,22,-66,3,-68,-36,-17,12,-30,0,-2,-25,-18,19,28,36,-37,9,-33,0,-18,-15,-2,21,20,9,59,32,-26,-12,-17,0,-50,-49,-11,-32,4,-33,17,76,46,2,2,-8,11,61,38,-25,-65,-32,-35,-31,2,-27,-42,20,46,86,17,25,21,-19,-19,14,27,33,8,17,-29,-11,23,-12,-16,-5,15,47,-27,35,-3,-3,-63,22,-7,6,12,-24,-7,-7,-31,75,87,29,-11,-39,52,36,-35,14,19,28,1,-3,23,-1,39,31,4,12,29,-35,-15,-1,17,13,56,-4,-22,-40,-34,-15,29,64,33,64,-13,-25,12,23,-43,37,0,25,-21,-15,25,-47,26,-5,25,-6,43,-53,0,-9,19,6,-41,-26,-27,-40,-7,-13,16,74,24,43,30,-67,60,-23,22,-80,-20,-30,15,-35,22,-23,32,4,-22,27,-6,-12,-62,-61,-4,-30,1,-13));
	end procedure get_input;
	
	procedure calculate_y(variable x_1D : in x_array_1D;
							variable w_2D : in w_array_2D;
							variable y_1D : out y_array_1D) IS
		
		variable accumulator : integer := 0;
		begin
			for i in 0 to 15 loop
				accumulator := 0;
				for j in 0 to 1023 loop
					accumulator := accumulator + w_2D(i,j)*x_1D(j);
				end loop;
				y_1D(i) := accumulator;
			end loop;
	end procedure calculate_y;

	procedure distance(variable y_1D : in y_array_1D;
						 variable yp_2D : in yp_array_2D;
						 variable index : out integer;
						 variable minNorm : out integer) IS
		variable dist : integer :=0;
		variable temp : integer :=0;
		variable minDist : integer := 99999999;
		begin
			index := -1;
			for i in 0 to 149 loop
				dist := 0;
				for j in 0 to 15 loop
					temp := yp_2D(i,j) - y_1D(j);
					if temp < 0 then
						dist := dist - temp;
					else
						dist := dist + temp;
					end if;
				end loop;
				
				if dist < minDist then
					minNorm := dist;
					minDist := dist;
					index := i;
				--else
					--minNorm := minNorm;
					--index := index;
				end if;
				
			end loop;
	end procedure distance;
			
end package body;
