--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   23:15:51 11/24/2016
-- Design Name:   
-- Module Name:   E:/14.7/ISE_DS/files/FaceRecoViaPCNN/tb_controlUnit.vhd
-- Project Name:  FaceRecoViaPCNN
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: ControlUnit
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY tb_controlUnit IS
END tb_controlUnit;
 
ARCHITECTURE behavior OF tb_controlUnit IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT ControlUnit
    PORT(
         clk : IN  std_logic;
         out_index : OUT  integer;
         slider : IN  integer;
         out_minNorm : OUT  integer
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal slider : integer := 0;

 	--Outputs
   signal out_index : integer;
   signal out_minNorm : integer;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: ControlUnit PORT MAP (
          clk => clk,
          out_index => out_index,
          slider => slider,
          out_minNorm => out_minNorm
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
		
		slider <= 0;
		wait for 50 ns;
		slider <= 1;
		wait for 50 ns;
		slider <= 2;
		wait for 50 ns;
		slider <= 3;
		wait for 50 ns;
		slider <= 4;
		wait for 50 ns;
		slider <= 5;
		wait for 50 ns;
		slider <= 6;
		wait for 50 ns;
		slider <= 7;
		wait for 50 ns;
		slider <= 8;
		wait for 50 ns;
		slider <= 9;
		wait for 50 ns;
		slider <= 10;
		wait for 50 ns;
		slider <= 11;
		wait for 50 ns;
		slider <= 12;
		wait for 50 ns;
		slider <= 13;
		wait for 50 ns;
		slider <= 14;
		wait for 50 ns;
		slider <= 15;
      wait for 100 ns;	

      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
